//File name  :    osmlgd_top.v
//Author     :    xiaocuicui
//Time       :    2022/05/21 14:10:24
//Version    :    V1.0
//Abstract   :        


`timescale 1ns/1ps

module osmlgd_top(clk,rst,work,
                  tx,
                  free, deout, valid);

//Define parameters:
parameter iteration = 10;
parameter rigth_formular = 0;

parameter init = 'd0;
parameter getin = 'd1;
parameter dot = 'd2;
parameter judge = 'd3;
parameter check = 'd4;
parameter compare = 'd5;
parameter update = 'd6;
parameter decode = 'd7;

//Define pins:
input clk;
input rst;
input work;
input [255:0] tx;
output wire free;
output wire [255:0] deout;
output wire valid;

//Define signals:
reg [2:0] state;

reg [255:0] Harray [127:0];
reg [255:0] tx_buffer;
reg [255:0] dotarray [127:0];
reg [127:0] form_array;
reg [7:0] check_cnt [255:0];
reg [7:0] wrong_cnt [255:0];
reg [255:0] update_buffer;
reg [3:0] iter_cnt;
reg free_flag, valid_flag, iter_flag;
reg [255:0] deout_reg;

assign free = free_flag;
assign valid = valid_flag;
assign deout = deout_reg;

//Instance

wire [8:0] row_sum_0, row_sum_1, row_sum_2, row_sum_3, row_sum_4, row_sum_5, row_sum_6, row_sum_7, 
           row_sum_8, row_sum_9, row_sum_10, row_sum_11, row_sum_12, row_sum_13, row_sum_14, row_sum_15, 
           row_sum_16, row_sum_17, row_sum_18, row_sum_19, row_sum_20, row_sum_21, row_sum_22, row_sum_23, 
           row_sum_24, row_sum_25, row_sum_26, row_sum_27, row_sum_28, row_sum_29, row_sum_30, row_sum_31, 
           row_sum_32, row_sum_33, row_sum_34, row_sum_35, row_sum_36, row_sum_37, row_sum_38, row_sum_39, 
           row_sum_40, row_sum_41, row_sum_42, row_sum_43, row_sum_44, row_sum_45, row_sum_46, row_sum_47, 
           row_sum_48, row_sum_49, row_sum_50, row_sum_51, row_sum_52, row_sum_53, row_sum_54, row_sum_55, 
           row_sum_56, row_sum_57, row_sum_58, row_sum_59, row_sum_60, row_sum_61, row_sum_62, row_sum_63, 
           row_sum_64, row_sum_65, row_sum_66, row_sum_67, row_sum_68, row_sum_69, row_sum_70, row_sum_71, 
           row_sum_72, row_sum_73, row_sum_74, row_sum_75, row_sum_76, row_sum_77, row_sum_78, row_sum_79, 
           row_sum_80, row_sum_81, row_sum_82, row_sum_83, row_sum_84, row_sum_85, row_sum_86, row_sum_87, 
           row_sum_88, row_sum_89, row_sum_90, row_sum_91, row_sum_92, row_sum_93, row_sum_94, row_sum_95, 
           row_sum_96, row_sum_97, row_sum_98, row_sum_99, row_sum_100, row_sum_101, row_sum_102, row_sum_103, 
           row_sum_104, row_sum_105, row_sum_106, row_sum_107, row_sum_108, row_sum_109, row_sum_110, row_sum_111, 
           row_sum_112, row_sum_113, row_sum_114, row_sum_115, row_sum_116, row_sum_117, row_sum_118, row_sum_119, 
           row_sum_120, row_sum_121, row_sum_122, row_sum_123, row_sum_124, row_sum_125, row_sum_126, row_sum_127;

wire [127:0] row_sum_lastbit;

assign row_sum_lastbit = {row_sum_0[0], row_sum_1[0], row_sum_2[0], row_sum_3[0], row_sum_4[0], row_sum_5[0], row_sum_6[0], row_sum_7[0], 
                          row_sum_8[0], row_sum_9[0], row_sum_10[0], row_sum_11[0], row_sum_12[0], row_sum_13[0], row_sum_14[0], row_sum_15[0], 
                          row_sum_16[0], row_sum_17[0], row_sum_18[0], row_sum_19[0], row_sum_20[0], row_sum_21[0], row_sum_22[0], row_sum_23[0], 
                          row_sum_24[0], row_sum_25[0], row_sum_26[0], row_sum_27[0], row_sum_28[0], row_sum_29[0], row_sum_30[0], row_sum_31[0], 
                          row_sum_32[0], row_sum_33[0], row_sum_34[0], row_sum_35[0], row_sum_36[0], row_sum_37[0], row_sum_38[0], row_sum_39[0], 
                          row_sum_40[0], row_sum_41[0], row_sum_42[0], row_sum_43[0], row_sum_44[0], row_sum_45[0], row_sum_46[0], row_sum_47[0], 
                          row_sum_48[0], row_sum_49[0], row_sum_50[0], row_sum_51[0], row_sum_52[0], row_sum_53[0], row_sum_54[0], row_sum_55[0], 
                          row_sum_56[0], row_sum_57[0], row_sum_58[0], row_sum_59[0], row_sum_60[0], row_sum_61[0], row_sum_62[0], row_sum_63[0], 
                          row_sum_64[0], row_sum_65[0], row_sum_66[0], row_sum_67[0], row_sum_68[0], row_sum_69[0], row_sum_70[0], row_sum_71[0], 
                          row_sum_72[0], row_sum_73[0], row_sum_74[0], row_sum_75[0], row_sum_76[0], row_sum_77[0], row_sum_78[0], row_sum_79[0], 
                          row_sum_80[0], row_sum_81[0], row_sum_82[0], row_sum_83[0], row_sum_84[0], row_sum_85[0], row_sum_86[0], row_sum_87[0], 
                          row_sum_88[0], row_sum_89[0], row_sum_90[0], row_sum_91[0], row_sum_92[0], row_sum_93[0], row_sum_94[0], row_sum_95[0], 
                          row_sum_96[0], row_sum_97[0], row_sum_98[0], row_sum_99[0], row_sum_100[0], row_sum_101[0], row_sum_102[0], row_sum_103[0], 
                          row_sum_104[0], row_sum_105[0], row_sum_106[0], row_sum_107[0], row_sum_108[0], row_sum_109[0], row_sum_110[0], row_sum_111[0], 
                          row_sum_112[0], row_sum_113[0], row_sum_114[0], row_sum_115[0], row_sum_116[0], row_sum_117[0], row_sum_118[0], row_sum_119[0], 
                          row_sum_120[0], row_sum_121[0], row_sum_122[0], row_sum_123[0], row_sum_124[0], row_sum_125[0], row_sum_126[0], row_sum_127[0]};


bitsadder_256 f_check_0(dotarray[0], row_sum_0);
bitsadder_256 f_check_1(dotarray[1], row_sum_1);
bitsadder_256 f_check_2(dotarray[2], row_sum_2);
bitsadder_256 f_check_3(dotarray[3], row_sum_3);
bitsadder_256 f_check_4(dotarray[4], row_sum_4);
bitsadder_256 f_check_5(dotarray[5], row_sum_5);
bitsadder_256 f_check_6(dotarray[6], row_sum_6);
bitsadder_256 f_check_7(dotarray[7], row_sum_7);
bitsadder_256 f_check_8(dotarray[8], row_sum_8);
bitsadder_256 f_check_9(dotarray[9], row_sum_9);
bitsadder_256 f_check_10(dotarray[10], row_sum_10);
bitsadder_256 f_check_11(dotarray[11], row_sum_11);
bitsadder_256 f_check_12(dotarray[12], row_sum_12);
bitsadder_256 f_check_13(dotarray[13], row_sum_13);
bitsadder_256 f_check_14(dotarray[14], row_sum_14);
bitsadder_256 f_check_15(dotarray[15], row_sum_15);
bitsadder_256 f_check_16(dotarray[16], row_sum_16);
bitsadder_256 f_check_17(dotarray[17], row_sum_17);
bitsadder_256 f_check_18(dotarray[18], row_sum_18);
bitsadder_256 f_check_19(dotarray[19], row_sum_19);
bitsadder_256 f_check_20(dotarray[20], row_sum_20);
bitsadder_256 f_check_21(dotarray[21], row_sum_21);
bitsadder_256 f_check_22(dotarray[22], row_sum_22);
bitsadder_256 f_check_23(dotarray[23], row_sum_23);
bitsadder_256 f_check_24(dotarray[24], row_sum_24);
bitsadder_256 f_check_25(dotarray[25], row_sum_25);
bitsadder_256 f_check_26(dotarray[26], row_sum_26);
bitsadder_256 f_check_27(dotarray[27], row_sum_27);
bitsadder_256 f_check_28(dotarray[28], row_sum_28);
bitsadder_256 f_check_29(dotarray[29], row_sum_29);
bitsadder_256 f_check_30(dotarray[30], row_sum_30);
bitsadder_256 f_check_31(dotarray[31], row_sum_31);
bitsadder_256 f_check_32(dotarray[32], row_sum_32);
bitsadder_256 f_check_33(dotarray[33], row_sum_33);
bitsadder_256 f_check_34(dotarray[34], row_sum_34);
bitsadder_256 f_check_35(dotarray[35], row_sum_35);
bitsadder_256 f_check_36(dotarray[36], row_sum_36);
bitsadder_256 f_check_37(dotarray[37], row_sum_37);
bitsadder_256 f_check_38(dotarray[38], row_sum_38);
bitsadder_256 f_check_39(dotarray[39], row_sum_39);
bitsadder_256 f_check_40(dotarray[40], row_sum_40);
bitsadder_256 f_check_41(dotarray[41], row_sum_41);
bitsadder_256 f_check_42(dotarray[42], row_sum_42);
bitsadder_256 f_check_43(dotarray[43], row_sum_43);
bitsadder_256 f_check_44(dotarray[44], row_sum_44);
bitsadder_256 f_check_45(dotarray[45], row_sum_45);
bitsadder_256 f_check_46(dotarray[46], row_sum_46);
bitsadder_256 f_check_47(dotarray[47], row_sum_47);
bitsadder_256 f_check_48(dotarray[48], row_sum_48);
bitsadder_256 f_check_49(dotarray[49], row_sum_49);
bitsadder_256 f_check_50(dotarray[50], row_sum_50);
bitsadder_256 f_check_51(dotarray[51], row_sum_51);
bitsadder_256 f_check_52(dotarray[52], row_sum_52);
bitsadder_256 f_check_53(dotarray[53], row_sum_53);
bitsadder_256 f_check_54(dotarray[54], row_sum_54);
bitsadder_256 f_check_55(dotarray[55], row_sum_55);
bitsadder_256 f_check_56(dotarray[56], row_sum_56);
bitsadder_256 f_check_57(dotarray[57], row_sum_57);
bitsadder_256 f_check_58(dotarray[58], row_sum_58);
bitsadder_256 f_check_59(dotarray[59], row_sum_59);
bitsadder_256 f_check_60(dotarray[60], row_sum_60);
bitsadder_256 f_check_61(dotarray[61], row_sum_61);
bitsadder_256 f_check_62(dotarray[62], row_sum_62);
bitsadder_256 f_check_63(dotarray[63], row_sum_63);
bitsadder_256 f_check_64(dotarray[64], row_sum_64);
bitsadder_256 f_check_65(dotarray[65], row_sum_65);
bitsadder_256 f_check_66(dotarray[66], row_sum_66);
bitsadder_256 f_check_67(dotarray[67], row_sum_67);
bitsadder_256 f_check_68(dotarray[68], row_sum_68);
bitsadder_256 f_check_69(dotarray[69], row_sum_69);
bitsadder_256 f_check_70(dotarray[70], row_sum_70);
bitsadder_256 f_check_71(dotarray[71], row_sum_71);
bitsadder_256 f_check_72(dotarray[72], row_sum_72);
bitsadder_256 f_check_73(dotarray[73], row_sum_73);
bitsadder_256 f_check_74(dotarray[74], row_sum_74);
bitsadder_256 f_check_75(dotarray[75], row_sum_75);
bitsadder_256 f_check_76(dotarray[76], row_sum_76);
bitsadder_256 f_check_77(dotarray[77], row_sum_77);
bitsadder_256 f_check_78(dotarray[78], row_sum_78);
bitsadder_256 f_check_79(dotarray[79], row_sum_79);
bitsadder_256 f_check_80(dotarray[80], row_sum_80);
bitsadder_256 f_check_81(dotarray[81], row_sum_81);
bitsadder_256 f_check_82(dotarray[82], row_sum_82);
bitsadder_256 f_check_83(dotarray[83], row_sum_83);
bitsadder_256 f_check_84(dotarray[84], row_sum_84);
bitsadder_256 f_check_85(dotarray[85], row_sum_85);
bitsadder_256 f_check_86(dotarray[86], row_sum_86);
bitsadder_256 f_check_87(dotarray[87], row_sum_87);
bitsadder_256 f_check_88(dotarray[88], row_sum_88);
bitsadder_256 f_check_89(dotarray[89], row_sum_89);
bitsadder_256 f_check_90(dotarray[90], row_sum_90);
bitsadder_256 f_check_91(dotarray[91], row_sum_91);
bitsadder_256 f_check_92(dotarray[92], row_sum_92);
bitsadder_256 f_check_93(dotarray[93], row_sum_93);
bitsadder_256 f_check_94(dotarray[94], row_sum_94);
bitsadder_256 f_check_95(dotarray[95], row_sum_95);
bitsadder_256 f_check_96(dotarray[96], row_sum_96);
bitsadder_256 f_check_97(dotarray[97], row_sum_97);
bitsadder_256 f_check_98(dotarray[98], row_sum_98);
bitsadder_256 f_check_99(dotarray[99], row_sum_99);
bitsadder_256 f_check_100(dotarray[100], row_sum_100);
bitsadder_256 f_check_101(dotarray[101], row_sum_101);
bitsadder_256 f_check_102(dotarray[102], row_sum_102);
bitsadder_256 f_check_103(dotarray[103], row_sum_103);
bitsadder_256 f_check_104(dotarray[104], row_sum_104);
bitsadder_256 f_check_105(dotarray[105], row_sum_105);
bitsadder_256 f_check_106(dotarray[106], row_sum_106);
bitsadder_256 f_check_107(dotarray[107], row_sum_107);
bitsadder_256 f_check_108(dotarray[108], row_sum_108);
bitsadder_256 f_check_109(dotarray[109], row_sum_109);
bitsadder_256 f_check_110(dotarray[110], row_sum_110);
bitsadder_256 f_check_111(dotarray[111], row_sum_111);
bitsadder_256 f_check_112(dotarray[112], row_sum_112);
bitsadder_256 f_check_113(dotarray[113], row_sum_113);
bitsadder_256 f_check_114(dotarray[114], row_sum_114);
bitsadder_256 f_check_115(dotarray[115], row_sum_115);
bitsadder_256 f_check_116(dotarray[116], row_sum_116);
bitsadder_256 f_check_117(dotarray[117], row_sum_117);
bitsadder_256 f_check_118(dotarray[118], row_sum_118);
bitsadder_256 f_check_119(dotarray[119], row_sum_119);
bitsadder_256 f_check_120(dotarray[120], row_sum_120);
bitsadder_256 f_check_121(dotarray[121], row_sum_121);
bitsadder_256 f_check_122(dotarray[122], row_sum_122);
bitsadder_256 f_check_123(dotarray[123], row_sum_123);
bitsadder_256 f_check_124(dotarray[124], row_sum_124);
bitsadder_256 f_check_125(dotarray[125], row_sum_125);
bitsadder_256 f_check_126(dotarray[126], row_sum_126);
bitsadder_256 f_check_127(dotarray[127], row_sum_127);

wire [127:0] h_col_0, h_col_1, h_col_2, h_col_3, h_col_4, h_col_5, h_col_6, h_col_7, 
             h_col_8, h_col_9, h_col_10, h_col_11, h_col_12, h_col_13, h_col_14, h_col_15, 
             h_col_16, h_col_17, h_col_18, h_col_19, h_col_20, h_col_21, h_col_22, h_col_23, 
             h_col_24, h_col_25, h_col_26, h_col_27, h_col_28, h_col_29, h_col_30, h_col_31, 
             h_col_32, h_col_33, h_col_34, h_col_35, h_col_36, h_col_37, h_col_38, h_col_39, 
             h_col_40, h_col_41, h_col_42, h_col_43, h_col_44, h_col_45, h_col_46, h_col_47, 
             h_col_48, h_col_49, h_col_50, h_col_51, h_col_52, h_col_53, h_col_54, h_col_55, 
             h_col_56, h_col_57, h_col_58, h_col_59, h_col_60, h_col_61, h_col_62, h_col_63, 
             h_col_64, h_col_65, h_col_66, h_col_67, h_col_68, h_col_69, h_col_70, h_col_71, 
             h_col_72, h_col_73, h_col_74, h_col_75, h_col_76, h_col_77, h_col_78, h_col_79, 
             h_col_80, h_col_81, h_col_82, h_col_83, h_col_84, h_col_85, h_col_86, h_col_87, 
             h_col_88, h_col_89, h_col_90, h_col_91, h_col_92, h_col_93, h_col_94, h_col_95, 
             h_col_96, h_col_97, h_col_98, h_col_99, h_col_100, h_col_101, h_col_102, h_col_103, 
             h_col_104, h_col_105, h_col_106, h_col_107, h_col_108, h_col_109, h_col_110, h_col_111, 
             h_col_112, h_col_113, h_col_114, h_col_115, h_col_116, h_col_117, h_col_118, h_col_119, 
             h_col_120, h_col_121, h_col_122, h_col_123, h_col_124, h_col_125, h_col_126, h_col_127, 
             h_col_128, h_col_129, h_col_130, h_col_131, h_col_132, h_col_133, h_col_134, h_col_135, 
             h_col_136, h_col_137, h_col_138, h_col_139, h_col_140, h_col_141, h_col_142, h_col_143, 
             h_col_144, h_col_145, h_col_146, h_col_147, h_col_148, h_col_149, h_col_150, h_col_151, 
             h_col_152, h_col_153, h_col_154, h_col_155, h_col_156, h_col_157, h_col_158, h_col_159, 
             h_col_160, h_col_161, h_col_162, h_col_163, h_col_164, h_col_165, h_col_166, h_col_167, 
             h_col_168, h_col_169, h_col_170, h_col_171, h_col_172, h_col_173, h_col_174, h_col_175, 
             h_col_176, h_col_177, h_col_178, h_col_179, h_col_180, h_col_181, h_col_182, h_col_183, 
             h_col_184, h_col_185, h_col_186, h_col_187, h_col_188, h_col_189, h_col_190, h_col_191, 
             h_col_192, h_col_193, h_col_194, h_col_195, h_col_196, h_col_197, h_col_198, h_col_199, 
             h_col_200, h_col_201, h_col_202, h_col_203, h_col_204, h_col_205, h_col_206, h_col_207, 
             h_col_208, h_col_209, h_col_210, h_col_211, h_col_212, h_col_213, h_col_214, h_col_215, 
             h_col_216, h_col_217, h_col_218, h_col_219, h_col_220, h_col_221, h_col_222, h_col_223, 
             h_col_224, h_col_225, h_col_226, h_col_227, h_col_228, h_col_229, h_col_230, h_col_231, 
             h_col_232, h_col_233, h_col_234, h_col_235, h_col_236, h_col_237, h_col_238, h_col_239, 
             h_col_240, h_col_241, h_col_242, h_col_243, h_col_244, h_col_245, h_col_246, h_col_247, 
             h_col_248, h_col_249, h_col_250, h_col_251, h_col_252, h_col_253, h_col_254, h_col_255;

assign h_col_0 = {Harray[0][0], Harray[1][0], Harray[2][0], Harray[3][0], Harray[4][0], Harray[5][0], Harray[6][0], Harray[7][0], Harray[8][0], Harray[9][0], Harray[10][0], Harray[11][0], Harray[12][0], Harray[13][0], Harray[14][0], Harray[15][0], Harray[16][0], Harray[17][0], Harray[18][0], Harray[19][0], Harray[20][0], Harray[21][0], Harray[22][0], Harray[23][0], Harray[24][0], Harray[25][0], Harray[26][0], Harray[27][0], Harray[28][0], Harray[29][0], Harray[30][0], Harray[31][0], Harray[32][0], Harray[33][0], Harray[34][0], Harray[35][0], Harray[36][0], Harray[37][0], Harray[38][0], Harray[39][0], Harray[40][0], Harray[41][0], Harray[42][0], Harray[43][0], Harray[44][0], Harray[45][0], Harray[46][0], Harray[47][0], Harray[48][0], Harray[49][0], Harray[50][0], Harray[51][0], Harray[52][0], Harray[53][0], Harray[54][0], Harray[55][0], Harray[56][0], Harray[57][0], Harray[58][0], Harray[59][0], Harray[60][0], Harray[61][0], Harray[62][0], Harray[63][0], Harray[64][0], Harray[65][0], Harray[66][0], Harray[67][0], Harray[68][0], Harray[69][0], Harray[70][0], Harray[71][0], Harray[72][0], Harray[73][0], Harray[74][0], Harray[75][0], Harray[76][0], Harray[77][0], Harray[78][0], Harray[79][0], Harray[80][0], Harray[81][0], Harray[82][0], Harray[83][0], Harray[84][0], Harray[85][0], Harray[86][0], Harray[87][0], Harray[88][0], Harray[89][0], Harray[90][0], Harray[91][0], Harray[92][0], Harray[93][0], Harray[94][0], Harray[95][0], Harray[96][0], Harray[97][0], Harray[98][0], Harray[99][0], Harray[100][0], Harray[101][0], Harray[102][0], Harray[103][0], Harray[104][0], Harray[105][0], Harray[106][0], Harray[107][0], Harray[108][0], Harray[109][0], Harray[110][0], Harray[111][0], Harray[112][0], Harray[113][0], Harray[114][0], Harray[115][0], Harray[116][0], Harray[117][0], Harray[118][0], Harray[119][0], Harray[120][0], Harray[121][0], Harray[122][0], Harray[123][0], Harray[124][0], Harray[125][0], Harray[126][0], Harray[127][0]};
assign h_col_1 = {Harray[0][1], Harray[1][1], Harray[2][1], Harray[3][1], Harray[4][1], Harray[5][1], Harray[6][1], Harray[7][1], Harray[8][1], Harray[9][1], Harray[10][1], Harray[11][1], Harray[12][1], Harray[13][1], Harray[14][1], Harray[15][1], Harray[16][1], Harray[17][1], Harray[18][1], Harray[19][1], Harray[20][1], Harray[21][1], Harray[22][1], Harray[23][1], Harray[24][1], Harray[25][1], Harray[26][1], Harray[27][1], Harray[28][1], Harray[29][1], Harray[30][1], Harray[31][1], Harray[32][1], Harray[33][1], Harray[34][1], Harray[35][1], Harray[36][1], Harray[37][1], Harray[38][1], Harray[39][1], Harray[40][1], Harray[41][1], Harray[42][1], Harray[43][1], Harray[44][1], Harray[45][1], Harray[46][1], Harray[47][1], Harray[48][1], Harray[49][1], Harray[50][1], Harray[51][1], Harray[52][1], Harray[53][1], Harray[54][1], Harray[55][1], Harray[56][1], Harray[57][1], Harray[58][1], Harray[59][1], Harray[60][1], Harray[61][1], Harray[62][1], Harray[63][1], Harray[64][1], Harray[65][1], Harray[66][1], Harray[67][1], Harray[68][1], Harray[69][1], Harray[70][1], Harray[71][1], Harray[72][1], Harray[73][1], Harray[74][1], Harray[75][1], Harray[76][1], Harray[77][1], Harray[78][1], Harray[79][1], Harray[80][1], Harray[81][1], Harray[82][1], Harray[83][1], Harray[84][1], Harray[85][1], Harray[86][1], Harray[87][1], Harray[88][1], Harray[89][1], Harray[90][1], Harray[91][1], Harray[92][1], Harray[93][1], Harray[94][1], Harray[95][1], Harray[96][1], Harray[97][1], Harray[98][1], Harray[99][1], Harray[100][1], Harray[101][1], Harray[102][1], Harray[103][1], Harray[104][1], Harray[105][1], Harray[106][1], Harray[107][1], Harray[108][1], Harray[109][1], Harray[110][1], Harray[111][1], Harray[112][1], Harray[113][1], Harray[114][1], Harray[115][1], Harray[116][1], Harray[117][1], Harray[118][1], Harray[119][1], Harray[120][1], Harray[121][1], Harray[122][1], Harray[123][1], Harray[124][1], Harray[125][1], Harray[126][1], Harray[127][1]};
assign h_col_2 = {Harray[0][2], Harray[1][2], Harray[2][2], Harray[3][2], Harray[4][2], Harray[5][2], Harray[6][2], Harray[7][2], Harray[8][2], Harray[9][2], Harray[10][2], Harray[11][2], Harray[12][2], Harray[13][2], Harray[14][2], Harray[15][2], Harray[16][2], Harray[17][2], Harray[18][2], Harray[19][2], Harray[20][2], Harray[21][2], Harray[22][2], Harray[23][2], Harray[24][2], Harray[25][2], Harray[26][2], Harray[27][2], Harray[28][2], Harray[29][2], Harray[30][2], Harray[31][2], Harray[32][2], Harray[33][2], Harray[34][2], Harray[35][2], Harray[36][2], Harray[37][2], Harray[38][2], Harray[39][2], Harray[40][2], Harray[41][2], Harray[42][2], Harray[43][2], Harray[44][2], Harray[45][2], Harray[46][2], Harray[47][2], Harray[48][2], Harray[49][2], Harray[50][2], Harray[51][2], Harray[52][2], Harray[53][2], Harray[54][2], Harray[55][2], Harray[56][2], Harray[57][2], Harray[58][2], Harray[59][2], Harray[60][2], Harray[61][2], Harray[62][2], Harray[63][2], Harray[64][2], Harray[65][2], Harray[66][2], Harray[67][2], Harray[68][2], Harray[69][2], Harray[70][2], Harray[71][2], Harray[72][2], Harray[73][2], Harray[74][2], Harray[75][2], Harray[76][2], Harray[77][2], Harray[78][2], Harray[79][2], Harray[80][2], Harray[81][2], Harray[82][2], Harray[83][2], Harray[84][2], Harray[85][2], Harray[86][2], Harray[87][2], Harray[88][2], Harray[89][2], Harray[90][2], Harray[91][2], Harray[92][2], Harray[93][2], Harray[94][2], Harray[95][2], Harray[96][2], Harray[97][2], Harray[98][2], Harray[99][2], Harray[100][2], Harray[101][2], Harray[102][2], Harray[103][2], Harray[104][2], Harray[105][2], Harray[106][2], Harray[107][2], Harray[108][2], Harray[109][2], Harray[110][2], Harray[111][2], Harray[112][2], Harray[113][2], Harray[114][2], Harray[115][2], Harray[116][2], Harray[117][2], Harray[118][2], Harray[119][2], Harray[120][2], Harray[121][2], Harray[122][2], Harray[123][2], Harray[124][2], Harray[125][2], Harray[126][2], Harray[127][2]};
assign h_col_3 = {Harray[0][3], Harray[1][3], Harray[2][3], Harray[3][3], Harray[4][3], Harray[5][3], Harray[6][3], Harray[7][3], Harray[8][3], Harray[9][3], Harray[10][3], Harray[11][3], Harray[12][3], Harray[13][3], Harray[14][3], Harray[15][3], Harray[16][3], Harray[17][3], Harray[18][3], Harray[19][3], Harray[20][3], Harray[21][3], Harray[22][3], Harray[23][3], Harray[24][3], Harray[25][3], Harray[26][3], Harray[27][3], Harray[28][3], Harray[29][3], Harray[30][3], Harray[31][3], Harray[32][3], Harray[33][3], Harray[34][3], Harray[35][3], Harray[36][3], Harray[37][3], Harray[38][3], Harray[39][3], Harray[40][3], Harray[41][3], Harray[42][3], Harray[43][3], Harray[44][3], Harray[45][3], Harray[46][3], Harray[47][3], Harray[48][3], Harray[49][3], Harray[50][3], Harray[51][3], Harray[52][3], Harray[53][3], Harray[54][3], Harray[55][3], Harray[56][3], Harray[57][3], Harray[58][3], Harray[59][3], Harray[60][3], Harray[61][3], Harray[62][3], Harray[63][3], Harray[64][3], Harray[65][3], Harray[66][3], Harray[67][3], Harray[68][3], Harray[69][3], Harray[70][3], Harray[71][3], Harray[72][3], Harray[73][3], Harray[74][3], Harray[75][3], Harray[76][3], Harray[77][3], Harray[78][3], Harray[79][3], Harray[80][3], Harray[81][3], Harray[82][3], Harray[83][3], Harray[84][3], Harray[85][3], Harray[86][3], Harray[87][3], Harray[88][3], Harray[89][3], Harray[90][3], Harray[91][3], Harray[92][3], Harray[93][3], Harray[94][3], Harray[95][3], Harray[96][3], Harray[97][3], Harray[98][3], Harray[99][3], Harray[100][3], Harray[101][3], Harray[102][3], Harray[103][3], Harray[104][3], Harray[105][3], Harray[106][3], Harray[107][3], Harray[108][3], Harray[109][3], Harray[110][3], Harray[111][3], Harray[112][3], Harray[113][3], Harray[114][3], Harray[115][3], Harray[116][3], Harray[117][3], Harray[118][3], Harray[119][3], Harray[120][3], Harray[121][3], Harray[122][3], Harray[123][3], Harray[124][3], Harray[125][3], Harray[126][3], Harray[127][3]};
assign h_col_4 = {Harray[0][4], Harray[1][4], Harray[2][4], Harray[3][4], Harray[4][4], Harray[5][4], Harray[6][4], Harray[7][4], Harray[8][4], Harray[9][4], Harray[10][4], Harray[11][4], Harray[12][4], Harray[13][4], Harray[14][4], Harray[15][4], Harray[16][4], Harray[17][4], Harray[18][4], Harray[19][4], Harray[20][4], Harray[21][4], Harray[22][4], Harray[23][4], Harray[24][4], Harray[25][4], Harray[26][4], Harray[27][4], Harray[28][4], Harray[29][4], Harray[30][4], Harray[31][4], Harray[32][4], Harray[33][4], Harray[34][4], Harray[35][4], Harray[36][4], Harray[37][4], Harray[38][4], Harray[39][4], Harray[40][4], Harray[41][4], Harray[42][4], Harray[43][4], Harray[44][4], Harray[45][4], Harray[46][4], Harray[47][4], Harray[48][4], Harray[49][4], Harray[50][4], Harray[51][4], Harray[52][4], Harray[53][4], Harray[54][4], Harray[55][4], Harray[56][4], Harray[57][4], Harray[58][4], Harray[59][4], Harray[60][4], Harray[61][4], Harray[62][4], Harray[63][4], Harray[64][4], Harray[65][4], Harray[66][4], Harray[67][4], Harray[68][4], Harray[69][4], Harray[70][4], Harray[71][4], Harray[72][4], Harray[73][4], Harray[74][4], Harray[75][4], Harray[76][4], Harray[77][4], Harray[78][4], Harray[79][4], Harray[80][4], Harray[81][4], Harray[82][4], Harray[83][4], Harray[84][4], Harray[85][4], Harray[86][4], Harray[87][4], Harray[88][4], Harray[89][4], Harray[90][4], Harray[91][4], Harray[92][4], Harray[93][4], Harray[94][4], Harray[95][4], Harray[96][4], Harray[97][4], Harray[98][4], Harray[99][4], Harray[100][4], Harray[101][4], Harray[102][4], Harray[103][4], Harray[104][4], Harray[105][4], Harray[106][4], Harray[107][4], Harray[108][4], Harray[109][4], Harray[110][4], Harray[111][4], Harray[112][4], Harray[113][4], Harray[114][4], Harray[115][4], Harray[116][4], Harray[117][4], Harray[118][4], Harray[119][4], Harray[120][4], Harray[121][4], Harray[122][4], Harray[123][4], Harray[124][4], Harray[125][4], Harray[126][4], Harray[127][4]};
assign h_col_5 = {Harray[0][5], Harray[1][5], Harray[2][5], Harray[3][5], Harray[4][5], Harray[5][5], Harray[6][5], Harray[7][5], Harray[8][5], Harray[9][5], Harray[10][5], Harray[11][5], Harray[12][5], Harray[13][5], Harray[14][5], Harray[15][5], Harray[16][5], Harray[17][5], Harray[18][5], Harray[19][5], Harray[20][5], Harray[21][5], Harray[22][5], Harray[23][5], Harray[24][5], Harray[25][5], Harray[26][5], Harray[27][5], Harray[28][5], Harray[29][5], Harray[30][5], Harray[31][5], Harray[32][5], Harray[33][5], Harray[34][5], Harray[35][5], Harray[36][5], Harray[37][5], Harray[38][5], Harray[39][5], Harray[40][5], Harray[41][5], Harray[42][5], Harray[43][5], Harray[44][5], Harray[45][5], Harray[46][5], Harray[47][5], Harray[48][5], Harray[49][5], Harray[50][5], Harray[51][5], Harray[52][5], Harray[53][5], Harray[54][5], Harray[55][5], Harray[56][5], Harray[57][5], Harray[58][5], Harray[59][5], Harray[60][5], Harray[61][5], Harray[62][5], Harray[63][5], Harray[64][5], Harray[65][5], Harray[66][5], Harray[67][5], Harray[68][5], Harray[69][5], Harray[70][5], Harray[71][5], Harray[72][5], Harray[73][5], Harray[74][5], Harray[75][5], Harray[76][5], Harray[77][5], Harray[78][5], Harray[79][5], Harray[80][5], Harray[81][5], Harray[82][5], Harray[83][5], Harray[84][5], Harray[85][5], Harray[86][5], Harray[87][5], Harray[88][5], Harray[89][5], Harray[90][5], Harray[91][5], Harray[92][5], Harray[93][5], Harray[94][5], Harray[95][5], Harray[96][5], Harray[97][5], Harray[98][5], Harray[99][5], Harray[100][5], Harray[101][5], Harray[102][5], Harray[103][5], Harray[104][5], Harray[105][5], Harray[106][5], Harray[107][5], Harray[108][5], Harray[109][5], Harray[110][5], Harray[111][5], Harray[112][5], Harray[113][5], Harray[114][5], Harray[115][5], Harray[116][5], Harray[117][5], Harray[118][5], Harray[119][5], Harray[120][5], Harray[121][5], Harray[122][5], Harray[123][5], Harray[124][5], Harray[125][5], Harray[126][5], Harray[127][5]};
assign h_col_6 = {Harray[0][6], Harray[1][6], Harray[2][6], Harray[3][6], Harray[4][6], Harray[5][6], Harray[6][6], Harray[7][6], Harray[8][6], Harray[9][6], Harray[10][6], Harray[11][6], Harray[12][6], Harray[13][6], Harray[14][6], Harray[15][6], Harray[16][6], Harray[17][6], Harray[18][6], Harray[19][6], Harray[20][6], Harray[21][6], Harray[22][6], Harray[23][6], Harray[24][6], Harray[25][6], Harray[26][6], Harray[27][6], Harray[28][6], Harray[29][6], Harray[30][6], Harray[31][6], Harray[32][6], Harray[33][6], Harray[34][6], Harray[35][6], Harray[36][6], Harray[37][6], Harray[38][6], Harray[39][6], Harray[40][6], Harray[41][6], Harray[42][6], Harray[43][6], Harray[44][6], Harray[45][6], Harray[46][6], Harray[47][6], Harray[48][6], Harray[49][6], Harray[50][6], Harray[51][6], Harray[52][6], Harray[53][6], Harray[54][6], Harray[55][6], Harray[56][6], Harray[57][6], Harray[58][6], Harray[59][6], Harray[60][6], Harray[61][6], Harray[62][6], Harray[63][6], Harray[64][6], Harray[65][6], Harray[66][6], Harray[67][6], Harray[68][6], Harray[69][6], Harray[70][6], Harray[71][6], Harray[72][6], Harray[73][6], Harray[74][6], Harray[75][6], Harray[76][6], Harray[77][6], Harray[78][6], Harray[79][6], Harray[80][6], Harray[81][6], Harray[82][6], Harray[83][6], Harray[84][6], Harray[85][6], Harray[86][6], Harray[87][6], Harray[88][6], Harray[89][6], Harray[90][6], Harray[91][6], Harray[92][6], Harray[93][6], Harray[94][6], Harray[95][6], Harray[96][6], Harray[97][6], Harray[98][6], Harray[99][6], Harray[100][6], Harray[101][6], Harray[102][6], Harray[103][6], Harray[104][6], Harray[105][6], Harray[106][6], Harray[107][6], Harray[108][6], Harray[109][6], Harray[110][6], Harray[111][6], Harray[112][6], Harray[113][6], Harray[114][6], Harray[115][6], Harray[116][6], Harray[117][6], Harray[118][6], Harray[119][6], Harray[120][6], Harray[121][6], Harray[122][6], Harray[123][6], Harray[124][6], Harray[125][6], Harray[126][6], Harray[127][6]};
assign h_col_7 = {Harray[0][7], Harray[1][7], Harray[2][7], Harray[3][7], Harray[4][7], Harray[5][7], Harray[6][7], Harray[7][7], Harray[8][7], Harray[9][7], Harray[10][7], Harray[11][7], Harray[12][7], Harray[13][7], Harray[14][7], Harray[15][7], Harray[16][7], Harray[17][7], Harray[18][7], Harray[19][7], Harray[20][7], Harray[21][7], Harray[22][7], Harray[23][7], Harray[24][7], Harray[25][7], Harray[26][7], Harray[27][7], Harray[28][7], Harray[29][7], Harray[30][7], Harray[31][7], Harray[32][7], Harray[33][7], Harray[34][7], Harray[35][7], Harray[36][7], Harray[37][7], Harray[38][7], Harray[39][7], Harray[40][7], Harray[41][7], Harray[42][7], Harray[43][7], Harray[44][7], Harray[45][7], Harray[46][7], Harray[47][7], Harray[48][7], Harray[49][7], Harray[50][7], Harray[51][7], Harray[52][7], Harray[53][7], Harray[54][7], Harray[55][7], Harray[56][7], Harray[57][7], Harray[58][7], Harray[59][7], Harray[60][7], Harray[61][7], Harray[62][7], Harray[63][7], Harray[64][7], Harray[65][7], Harray[66][7], Harray[67][7], Harray[68][7], Harray[69][7], Harray[70][7], Harray[71][7], Harray[72][7], Harray[73][7], Harray[74][7], Harray[75][7], Harray[76][7], Harray[77][7], Harray[78][7], Harray[79][7], Harray[80][7], Harray[81][7], Harray[82][7], Harray[83][7], Harray[84][7], Harray[85][7], Harray[86][7], Harray[87][7], Harray[88][7], Harray[89][7], Harray[90][7], Harray[91][7], Harray[92][7], Harray[93][7], Harray[94][7], Harray[95][7], Harray[96][7], Harray[97][7], Harray[98][7], Harray[99][7], Harray[100][7], Harray[101][7], Harray[102][7], Harray[103][7], Harray[104][7], Harray[105][7], Harray[106][7], Harray[107][7], Harray[108][7], Harray[109][7], Harray[110][7], Harray[111][7], Harray[112][7], Harray[113][7], Harray[114][7], Harray[115][7], Harray[116][7], Harray[117][7], Harray[118][7], Harray[119][7], Harray[120][7], Harray[121][7], Harray[122][7], Harray[123][7], Harray[124][7], Harray[125][7], Harray[126][7], Harray[127][7]};
assign h_col_8 = {Harray[0][8], Harray[1][8], Harray[2][8], Harray[3][8], Harray[4][8], Harray[5][8], Harray[6][8], Harray[7][8], Harray[8][8], Harray[9][8], Harray[10][8], Harray[11][8], Harray[12][8], Harray[13][8], Harray[14][8], Harray[15][8], Harray[16][8], Harray[17][8], Harray[18][8], Harray[19][8], Harray[20][8], Harray[21][8], Harray[22][8], Harray[23][8], Harray[24][8], Harray[25][8], Harray[26][8], Harray[27][8], Harray[28][8], Harray[29][8], Harray[30][8], Harray[31][8], Harray[32][8], Harray[33][8], Harray[34][8], Harray[35][8], Harray[36][8], Harray[37][8], Harray[38][8], Harray[39][8], Harray[40][8], Harray[41][8], Harray[42][8], Harray[43][8], Harray[44][8], Harray[45][8], Harray[46][8], Harray[47][8], Harray[48][8], Harray[49][8], Harray[50][8], Harray[51][8], Harray[52][8], Harray[53][8], Harray[54][8], Harray[55][8], Harray[56][8], Harray[57][8], Harray[58][8], Harray[59][8], Harray[60][8], Harray[61][8], Harray[62][8], Harray[63][8], Harray[64][8], Harray[65][8], Harray[66][8], Harray[67][8], Harray[68][8], Harray[69][8], Harray[70][8], Harray[71][8], Harray[72][8], Harray[73][8], Harray[74][8], Harray[75][8], Harray[76][8], Harray[77][8], Harray[78][8], Harray[79][8], Harray[80][8], Harray[81][8], Harray[82][8], Harray[83][8], Harray[84][8], Harray[85][8], Harray[86][8], Harray[87][8], Harray[88][8], Harray[89][8], Harray[90][8], Harray[91][8], Harray[92][8], Harray[93][8], Harray[94][8], Harray[95][8], Harray[96][8], Harray[97][8], Harray[98][8], Harray[99][8], Harray[100][8], Harray[101][8], Harray[102][8], Harray[103][8], Harray[104][8], Harray[105][8], Harray[106][8], Harray[107][8], Harray[108][8], Harray[109][8], Harray[110][8], Harray[111][8], Harray[112][8], Harray[113][8], Harray[114][8], Harray[115][8], Harray[116][8], Harray[117][8], Harray[118][8], Harray[119][8], Harray[120][8], Harray[121][8], Harray[122][8], Harray[123][8], Harray[124][8], Harray[125][8], Harray[126][8], Harray[127][8]};
assign h_col_9 = {Harray[0][9], Harray[1][9], Harray[2][9], Harray[3][9], Harray[4][9], Harray[5][9], Harray[6][9], Harray[7][9], Harray[8][9], Harray[9][9], Harray[10][9], Harray[11][9], Harray[12][9], Harray[13][9], Harray[14][9], Harray[15][9], Harray[16][9], Harray[17][9], Harray[18][9], Harray[19][9], Harray[20][9], Harray[21][9], Harray[22][9], Harray[23][9], Harray[24][9], Harray[25][9], Harray[26][9], Harray[27][9], Harray[28][9], Harray[29][9], Harray[30][9], Harray[31][9], Harray[32][9], Harray[33][9], Harray[34][9], Harray[35][9], Harray[36][9], Harray[37][9], Harray[38][9], Harray[39][9], Harray[40][9], Harray[41][9], Harray[42][9], Harray[43][9], Harray[44][9], Harray[45][9], Harray[46][9], Harray[47][9], Harray[48][9], Harray[49][9], Harray[50][9], Harray[51][9], Harray[52][9], Harray[53][9], Harray[54][9], Harray[55][9], Harray[56][9], Harray[57][9], Harray[58][9], Harray[59][9], Harray[60][9], Harray[61][9], Harray[62][9], Harray[63][9], Harray[64][9], Harray[65][9], Harray[66][9], Harray[67][9], Harray[68][9], Harray[69][9], Harray[70][9], Harray[71][9], Harray[72][9], Harray[73][9], Harray[74][9], Harray[75][9], Harray[76][9], Harray[77][9], Harray[78][9], Harray[79][9], Harray[80][9], Harray[81][9], Harray[82][9], Harray[83][9], Harray[84][9], Harray[85][9], Harray[86][9], Harray[87][9], Harray[88][9], Harray[89][9], Harray[90][9], Harray[91][9], Harray[92][9], Harray[93][9], Harray[94][9], Harray[95][9], Harray[96][9], Harray[97][9], Harray[98][9], Harray[99][9], Harray[100][9], Harray[101][9], Harray[102][9], Harray[103][9], Harray[104][9], Harray[105][9], Harray[106][9], Harray[107][9], Harray[108][9], Harray[109][9], Harray[110][9], Harray[111][9], Harray[112][9], Harray[113][9], Harray[114][9], Harray[115][9], Harray[116][9], Harray[117][9], Harray[118][9], Harray[119][9], Harray[120][9], Harray[121][9], Harray[122][9], Harray[123][9], Harray[124][9], Harray[125][9], Harray[126][9], Harray[127][9]};
assign h_col_10 = {Harray[0][10], Harray[1][10], Harray[2][10], Harray[3][10], Harray[4][10], Harray[5][10], Harray[6][10], Harray[7][10], Harray[8][10], Harray[9][10], Harray[10][10], Harray[11][10], Harray[12][10], Harray[13][10], Harray[14][10], Harray[15][10], Harray[16][10], Harray[17][10], Harray[18][10], Harray[19][10], Harray[20][10], Harray[21][10], Harray[22][10], Harray[23][10], Harray[24][10], Harray[25][10], Harray[26][10], Harray[27][10], Harray[28][10], Harray[29][10], Harray[30][10], Harray[31][10], Harray[32][10], Harray[33][10], Harray[34][10], Harray[35][10], Harray[36][10], Harray[37][10], Harray[38][10], Harray[39][10], Harray[40][10], Harray[41][10], Harray[42][10], Harray[43][10], Harray[44][10], Harray[45][10], Harray[46][10], Harray[47][10], Harray[48][10], Harray[49][10], Harray[50][10], Harray[51][10], Harray[52][10], Harray[53][10], Harray[54][10], Harray[55][10], Harray[56][10], Harray[57][10], Harray[58][10], Harray[59][10], Harray[60][10], Harray[61][10], Harray[62][10], Harray[63][10], Harray[64][10], Harray[65][10], Harray[66][10], Harray[67][10], Harray[68][10], Harray[69][10], Harray[70][10], Harray[71][10], Harray[72][10], Harray[73][10], Harray[74][10], Harray[75][10], Harray[76][10], Harray[77][10], Harray[78][10], Harray[79][10], Harray[80][10], Harray[81][10], Harray[82][10], Harray[83][10], Harray[84][10], Harray[85][10], Harray[86][10], Harray[87][10], Harray[88][10], Harray[89][10], Harray[90][10], Harray[91][10], Harray[92][10], Harray[93][10], Harray[94][10], Harray[95][10], Harray[96][10], Harray[97][10], Harray[98][10], Harray[99][10], Harray[100][10], Harray[101][10], Harray[102][10], Harray[103][10], Harray[104][10], Harray[105][10], Harray[106][10], Harray[107][10], Harray[108][10], Harray[109][10], Harray[110][10], Harray[111][10], Harray[112][10], Harray[113][10], Harray[114][10], Harray[115][10], Harray[116][10], Harray[117][10], Harray[118][10], Harray[119][10], Harray[120][10], Harray[121][10], Harray[122][10], Harray[123][10], Harray[124][10], Harray[125][10], Harray[126][10], Harray[127][10]};
assign h_col_11 = {Harray[0][11], Harray[1][11], Harray[2][11], Harray[3][11], Harray[4][11], Harray[5][11], Harray[6][11], Harray[7][11], Harray[8][11], Harray[9][11], Harray[10][11], Harray[11][11], Harray[12][11], Harray[13][11], Harray[14][11], Harray[15][11], Harray[16][11], Harray[17][11], Harray[18][11], Harray[19][11], Harray[20][11], Harray[21][11], Harray[22][11], Harray[23][11], Harray[24][11], Harray[25][11], Harray[26][11], Harray[27][11], Harray[28][11], Harray[29][11], Harray[30][11], Harray[31][11], Harray[32][11], Harray[33][11], Harray[34][11], Harray[35][11], Harray[36][11], Harray[37][11], Harray[38][11], Harray[39][11], Harray[40][11], Harray[41][11], Harray[42][11], Harray[43][11], Harray[44][11], Harray[45][11], Harray[46][11], Harray[47][11], Harray[48][11], Harray[49][11], Harray[50][11], Harray[51][11], Harray[52][11], Harray[53][11], Harray[54][11], Harray[55][11], Harray[56][11], Harray[57][11], Harray[58][11], Harray[59][11], Harray[60][11], Harray[61][11], Harray[62][11], Harray[63][11], Harray[64][11], Harray[65][11], Harray[66][11], Harray[67][11], Harray[68][11], Harray[69][11], Harray[70][11], Harray[71][11], Harray[72][11], Harray[73][11], Harray[74][11], Harray[75][11], Harray[76][11], Harray[77][11], Harray[78][11], Harray[79][11], Harray[80][11], Harray[81][11], Harray[82][11], Harray[83][11], Harray[84][11], Harray[85][11], Harray[86][11], Harray[87][11], Harray[88][11], Harray[89][11], Harray[90][11], Harray[91][11], Harray[92][11], Harray[93][11], Harray[94][11], Harray[95][11], Harray[96][11], Harray[97][11], Harray[98][11], Harray[99][11], Harray[100][11], Harray[101][11], Harray[102][11], Harray[103][11], Harray[104][11], Harray[105][11], Harray[106][11], Harray[107][11], Harray[108][11], Harray[109][11], Harray[110][11], Harray[111][11], Harray[112][11], Harray[113][11], Harray[114][11], Harray[115][11], Harray[116][11], Harray[117][11], Harray[118][11], Harray[119][11], Harray[120][11], Harray[121][11], Harray[122][11], Harray[123][11], Harray[124][11], Harray[125][11], Harray[126][11], Harray[127][11]};
assign h_col_12 = {Harray[0][12], Harray[1][12], Harray[2][12], Harray[3][12], Harray[4][12], Harray[5][12], Harray[6][12], Harray[7][12], Harray[8][12], Harray[9][12], Harray[10][12], Harray[11][12], Harray[12][12], Harray[13][12], Harray[14][12], Harray[15][12], Harray[16][12], Harray[17][12], Harray[18][12], Harray[19][12], Harray[20][12], Harray[21][12], Harray[22][12], Harray[23][12], Harray[24][12], Harray[25][12], Harray[26][12], Harray[27][12], Harray[28][12], Harray[29][12], Harray[30][12], Harray[31][12], Harray[32][12], Harray[33][12], Harray[34][12], Harray[35][12], Harray[36][12], Harray[37][12], Harray[38][12], Harray[39][12], Harray[40][12], Harray[41][12], Harray[42][12], Harray[43][12], Harray[44][12], Harray[45][12], Harray[46][12], Harray[47][12], Harray[48][12], Harray[49][12], Harray[50][12], Harray[51][12], Harray[52][12], Harray[53][12], Harray[54][12], Harray[55][12], Harray[56][12], Harray[57][12], Harray[58][12], Harray[59][12], Harray[60][12], Harray[61][12], Harray[62][12], Harray[63][12], Harray[64][12], Harray[65][12], Harray[66][12], Harray[67][12], Harray[68][12], Harray[69][12], Harray[70][12], Harray[71][12], Harray[72][12], Harray[73][12], Harray[74][12], Harray[75][12], Harray[76][12], Harray[77][12], Harray[78][12], Harray[79][12], Harray[80][12], Harray[81][12], Harray[82][12], Harray[83][12], Harray[84][12], Harray[85][12], Harray[86][12], Harray[87][12], Harray[88][12], Harray[89][12], Harray[90][12], Harray[91][12], Harray[92][12], Harray[93][12], Harray[94][12], Harray[95][12], Harray[96][12], Harray[97][12], Harray[98][12], Harray[99][12], Harray[100][12], Harray[101][12], Harray[102][12], Harray[103][12], Harray[104][12], Harray[105][12], Harray[106][12], Harray[107][12], Harray[108][12], Harray[109][12], Harray[110][12], Harray[111][12], Harray[112][12], Harray[113][12], Harray[114][12], Harray[115][12], Harray[116][12], Harray[117][12], Harray[118][12], Harray[119][12], Harray[120][12], Harray[121][12], Harray[122][12], Harray[123][12], Harray[124][12], Harray[125][12], Harray[126][12], Harray[127][12]};
assign h_col_13 = {Harray[0][13], Harray[1][13], Harray[2][13], Harray[3][13], Harray[4][13], Harray[5][13], Harray[6][13], Harray[7][13], Harray[8][13], Harray[9][13], Harray[10][13], Harray[11][13], Harray[12][13], Harray[13][13], Harray[14][13], Harray[15][13], Harray[16][13], Harray[17][13], Harray[18][13], Harray[19][13], Harray[20][13], Harray[21][13], Harray[22][13], Harray[23][13], Harray[24][13], Harray[25][13], Harray[26][13], Harray[27][13], Harray[28][13], Harray[29][13], Harray[30][13], Harray[31][13], Harray[32][13], Harray[33][13], Harray[34][13], Harray[35][13], Harray[36][13], Harray[37][13], Harray[38][13], Harray[39][13], Harray[40][13], Harray[41][13], Harray[42][13], Harray[43][13], Harray[44][13], Harray[45][13], Harray[46][13], Harray[47][13], Harray[48][13], Harray[49][13], Harray[50][13], Harray[51][13], Harray[52][13], Harray[53][13], Harray[54][13], Harray[55][13], Harray[56][13], Harray[57][13], Harray[58][13], Harray[59][13], Harray[60][13], Harray[61][13], Harray[62][13], Harray[63][13], Harray[64][13], Harray[65][13], Harray[66][13], Harray[67][13], Harray[68][13], Harray[69][13], Harray[70][13], Harray[71][13], Harray[72][13], Harray[73][13], Harray[74][13], Harray[75][13], Harray[76][13], Harray[77][13], Harray[78][13], Harray[79][13], Harray[80][13], Harray[81][13], Harray[82][13], Harray[83][13], Harray[84][13], Harray[85][13], Harray[86][13], Harray[87][13], Harray[88][13], Harray[89][13], Harray[90][13], Harray[91][13], Harray[92][13], Harray[93][13], Harray[94][13], Harray[95][13], Harray[96][13], Harray[97][13], Harray[98][13], Harray[99][13], Harray[100][13], Harray[101][13], Harray[102][13], Harray[103][13], Harray[104][13], Harray[105][13], Harray[106][13], Harray[107][13], Harray[108][13], Harray[109][13], Harray[110][13], Harray[111][13], Harray[112][13], Harray[113][13], Harray[114][13], Harray[115][13], Harray[116][13], Harray[117][13], Harray[118][13], Harray[119][13], Harray[120][13], Harray[121][13], Harray[122][13], Harray[123][13], Harray[124][13], Harray[125][13], Harray[126][13], Harray[127][13]};
assign h_col_14 = {Harray[0][14], Harray[1][14], Harray[2][14], Harray[3][14], Harray[4][14], Harray[5][14], Harray[6][14], Harray[7][14], Harray[8][14], Harray[9][14], Harray[10][14], Harray[11][14], Harray[12][14], Harray[13][14], Harray[14][14], Harray[15][14], Harray[16][14], Harray[17][14], Harray[18][14], Harray[19][14], Harray[20][14], Harray[21][14], Harray[22][14], Harray[23][14], Harray[24][14], Harray[25][14], Harray[26][14], Harray[27][14], Harray[28][14], Harray[29][14], Harray[30][14], Harray[31][14], Harray[32][14], Harray[33][14], Harray[34][14], Harray[35][14], Harray[36][14], Harray[37][14], Harray[38][14], Harray[39][14], Harray[40][14], Harray[41][14], Harray[42][14], Harray[43][14], Harray[44][14], Harray[45][14], Harray[46][14], Harray[47][14], Harray[48][14], Harray[49][14], Harray[50][14], Harray[51][14], Harray[52][14], Harray[53][14], Harray[54][14], Harray[55][14], Harray[56][14], Harray[57][14], Harray[58][14], Harray[59][14], Harray[60][14], Harray[61][14], Harray[62][14], Harray[63][14], Harray[64][14], Harray[65][14], Harray[66][14], Harray[67][14], Harray[68][14], Harray[69][14], Harray[70][14], Harray[71][14], Harray[72][14], Harray[73][14], Harray[74][14], Harray[75][14], Harray[76][14], Harray[77][14], Harray[78][14], Harray[79][14], Harray[80][14], Harray[81][14], Harray[82][14], Harray[83][14], Harray[84][14], Harray[85][14], Harray[86][14], Harray[87][14], Harray[88][14], Harray[89][14], Harray[90][14], Harray[91][14], Harray[92][14], Harray[93][14], Harray[94][14], Harray[95][14], Harray[96][14], Harray[97][14], Harray[98][14], Harray[99][14], Harray[100][14], Harray[101][14], Harray[102][14], Harray[103][14], Harray[104][14], Harray[105][14], Harray[106][14], Harray[107][14], Harray[108][14], Harray[109][14], Harray[110][14], Harray[111][14], Harray[112][14], Harray[113][14], Harray[114][14], Harray[115][14], Harray[116][14], Harray[117][14], Harray[118][14], Harray[119][14], Harray[120][14], Harray[121][14], Harray[122][14], Harray[123][14], Harray[124][14], Harray[125][14], Harray[126][14], Harray[127][14]};
assign h_col_15 = {Harray[0][15], Harray[1][15], Harray[2][15], Harray[3][15], Harray[4][15], Harray[5][15], Harray[6][15], Harray[7][15], Harray[8][15], Harray[9][15], Harray[10][15], Harray[11][15], Harray[12][15], Harray[13][15], Harray[14][15], Harray[15][15], Harray[16][15], Harray[17][15], Harray[18][15], Harray[19][15], Harray[20][15], Harray[21][15], Harray[22][15], Harray[23][15], Harray[24][15], Harray[25][15], Harray[26][15], Harray[27][15], Harray[28][15], Harray[29][15], Harray[30][15], Harray[31][15], Harray[32][15], Harray[33][15], Harray[34][15], Harray[35][15], Harray[36][15], Harray[37][15], Harray[38][15], Harray[39][15], Harray[40][15], Harray[41][15], Harray[42][15], Harray[43][15], Harray[44][15], Harray[45][15], Harray[46][15], Harray[47][15], Harray[48][15], Harray[49][15], Harray[50][15], Harray[51][15], Harray[52][15], Harray[53][15], Harray[54][15], Harray[55][15], Harray[56][15], Harray[57][15], Harray[58][15], Harray[59][15], Harray[60][15], Harray[61][15], Harray[62][15], Harray[63][15], Harray[64][15], Harray[65][15], Harray[66][15], Harray[67][15], Harray[68][15], Harray[69][15], Harray[70][15], Harray[71][15], Harray[72][15], Harray[73][15], Harray[74][15], Harray[75][15], Harray[76][15], Harray[77][15], Harray[78][15], Harray[79][15], Harray[80][15], Harray[81][15], Harray[82][15], Harray[83][15], Harray[84][15], Harray[85][15], Harray[86][15], Harray[87][15], Harray[88][15], Harray[89][15], Harray[90][15], Harray[91][15], Harray[92][15], Harray[93][15], Harray[94][15], Harray[95][15], Harray[96][15], Harray[97][15], Harray[98][15], Harray[99][15], Harray[100][15], Harray[101][15], Harray[102][15], Harray[103][15], Harray[104][15], Harray[105][15], Harray[106][15], Harray[107][15], Harray[108][15], Harray[109][15], Harray[110][15], Harray[111][15], Harray[112][15], Harray[113][15], Harray[114][15], Harray[115][15], Harray[116][15], Harray[117][15], Harray[118][15], Harray[119][15], Harray[120][15], Harray[121][15], Harray[122][15], Harray[123][15], Harray[124][15], Harray[125][15], Harray[126][15], Harray[127][15]};
assign h_col_16 = {Harray[0][16], Harray[1][16], Harray[2][16], Harray[3][16], Harray[4][16], Harray[5][16], Harray[6][16], Harray[7][16], Harray[8][16], Harray[9][16], Harray[10][16], Harray[11][16], Harray[12][16], Harray[13][16], Harray[14][16], Harray[15][16], Harray[16][16], Harray[17][16], Harray[18][16], Harray[19][16], Harray[20][16], Harray[21][16], Harray[22][16], Harray[23][16], Harray[24][16], Harray[25][16], Harray[26][16], Harray[27][16], Harray[28][16], Harray[29][16], Harray[30][16], Harray[31][16], Harray[32][16], Harray[33][16], Harray[34][16], Harray[35][16], Harray[36][16], Harray[37][16], Harray[38][16], Harray[39][16], Harray[40][16], Harray[41][16], Harray[42][16], Harray[43][16], Harray[44][16], Harray[45][16], Harray[46][16], Harray[47][16], Harray[48][16], Harray[49][16], Harray[50][16], Harray[51][16], Harray[52][16], Harray[53][16], Harray[54][16], Harray[55][16], Harray[56][16], Harray[57][16], Harray[58][16], Harray[59][16], Harray[60][16], Harray[61][16], Harray[62][16], Harray[63][16], Harray[64][16], Harray[65][16], Harray[66][16], Harray[67][16], Harray[68][16], Harray[69][16], Harray[70][16], Harray[71][16], Harray[72][16], Harray[73][16], Harray[74][16], Harray[75][16], Harray[76][16], Harray[77][16], Harray[78][16], Harray[79][16], Harray[80][16], Harray[81][16], Harray[82][16], Harray[83][16], Harray[84][16], Harray[85][16], Harray[86][16], Harray[87][16], Harray[88][16], Harray[89][16], Harray[90][16], Harray[91][16], Harray[92][16], Harray[93][16], Harray[94][16], Harray[95][16], Harray[96][16], Harray[97][16], Harray[98][16], Harray[99][16], Harray[100][16], Harray[101][16], Harray[102][16], Harray[103][16], Harray[104][16], Harray[105][16], Harray[106][16], Harray[107][16], Harray[108][16], Harray[109][16], Harray[110][16], Harray[111][16], Harray[112][16], Harray[113][16], Harray[114][16], Harray[115][16], Harray[116][16], Harray[117][16], Harray[118][16], Harray[119][16], Harray[120][16], Harray[121][16], Harray[122][16], Harray[123][16], Harray[124][16], Harray[125][16], Harray[126][16], Harray[127][16]};
assign h_col_17 = {Harray[0][17], Harray[1][17], Harray[2][17], Harray[3][17], Harray[4][17], Harray[5][17], Harray[6][17], Harray[7][17], Harray[8][17], Harray[9][17], Harray[10][17], Harray[11][17], Harray[12][17], Harray[13][17], Harray[14][17], Harray[15][17], Harray[16][17], Harray[17][17], Harray[18][17], Harray[19][17], Harray[20][17], Harray[21][17], Harray[22][17], Harray[23][17], Harray[24][17], Harray[25][17], Harray[26][17], Harray[27][17], Harray[28][17], Harray[29][17], Harray[30][17], Harray[31][17], Harray[32][17], Harray[33][17], Harray[34][17], Harray[35][17], Harray[36][17], Harray[37][17], Harray[38][17], Harray[39][17], Harray[40][17], Harray[41][17], Harray[42][17], Harray[43][17], Harray[44][17], Harray[45][17], Harray[46][17], Harray[47][17], Harray[48][17], Harray[49][17], Harray[50][17], Harray[51][17], Harray[52][17], Harray[53][17], Harray[54][17], Harray[55][17], Harray[56][17], Harray[57][17], Harray[58][17], Harray[59][17], Harray[60][17], Harray[61][17], Harray[62][17], Harray[63][17], Harray[64][17], Harray[65][17], Harray[66][17], Harray[67][17], Harray[68][17], Harray[69][17], Harray[70][17], Harray[71][17], Harray[72][17], Harray[73][17], Harray[74][17], Harray[75][17], Harray[76][17], Harray[77][17], Harray[78][17], Harray[79][17], Harray[80][17], Harray[81][17], Harray[82][17], Harray[83][17], Harray[84][17], Harray[85][17], Harray[86][17], Harray[87][17], Harray[88][17], Harray[89][17], Harray[90][17], Harray[91][17], Harray[92][17], Harray[93][17], Harray[94][17], Harray[95][17], Harray[96][17], Harray[97][17], Harray[98][17], Harray[99][17], Harray[100][17], Harray[101][17], Harray[102][17], Harray[103][17], Harray[104][17], Harray[105][17], Harray[106][17], Harray[107][17], Harray[108][17], Harray[109][17], Harray[110][17], Harray[111][17], Harray[112][17], Harray[113][17], Harray[114][17], Harray[115][17], Harray[116][17], Harray[117][17], Harray[118][17], Harray[119][17], Harray[120][17], Harray[121][17], Harray[122][17], Harray[123][17], Harray[124][17], Harray[125][17], Harray[126][17], Harray[127][17]};
assign h_col_18 = {Harray[0][18], Harray[1][18], Harray[2][18], Harray[3][18], Harray[4][18], Harray[5][18], Harray[6][18], Harray[7][18], Harray[8][18], Harray[9][18], Harray[10][18], Harray[11][18], Harray[12][18], Harray[13][18], Harray[14][18], Harray[15][18], Harray[16][18], Harray[17][18], Harray[18][18], Harray[19][18], Harray[20][18], Harray[21][18], Harray[22][18], Harray[23][18], Harray[24][18], Harray[25][18], Harray[26][18], Harray[27][18], Harray[28][18], Harray[29][18], Harray[30][18], Harray[31][18], Harray[32][18], Harray[33][18], Harray[34][18], Harray[35][18], Harray[36][18], Harray[37][18], Harray[38][18], Harray[39][18], Harray[40][18], Harray[41][18], Harray[42][18], Harray[43][18], Harray[44][18], Harray[45][18], Harray[46][18], Harray[47][18], Harray[48][18], Harray[49][18], Harray[50][18], Harray[51][18], Harray[52][18], Harray[53][18], Harray[54][18], Harray[55][18], Harray[56][18], Harray[57][18], Harray[58][18], Harray[59][18], Harray[60][18], Harray[61][18], Harray[62][18], Harray[63][18], Harray[64][18], Harray[65][18], Harray[66][18], Harray[67][18], Harray[68][18], Harray[69][18], Harray[70][18], Harray[71][18], Harray[72][18], Harray[73][18], Harray[74][18], Harray[75][18], Harray[76][18], Harray[77][18], Harray[78][18], Harray[79][18], Harray[80][18], Harray[81][18], Harray[82][18], Harray[83][18], Harray[84][18], Harray[85][18], Harray[86][18], Harray[87][18], Harray[88][18], Harray[89][18], Harray[90][18], Harray[91][18], Harray[92][18], Harray[93][18], Harray[94][18], Harray[95][18], Harray[96][18], Harray[97][18], Harray[98][18], Harray[99][18], Harray[100][18], Harray[101][18], Harray[102][18], Harray[103][18], Harray[104][18], Harray[105][18], Harray[106][18], Harray[107][18], Harray[108][18], Harray[109][18], Harray[110][18], Harray[111][18], Harray[112][18], Harray[113][18], Harray[114][18], Harray[115][18], Harray[116][18], Harray[117][18], Harray[118][18], Harray[119][18], Harray[120][18], Harray[121][18], Harray[122][18], Harray[123][18], Harray[124][18], Harray[125][18], Harray[126][18], Harray[127][18]};
assign h_col_19 = {Harray[0][19], Harray[1][19], Harray[2][19], Harray[3][19], Harray[4][19], Harray[5][19], Harray[6][19], Harray[7][19], Harray[8][19], Harray[9][19], Harray[10][19], Harray[11][19], Harray[12][19], Harray[13][19], Harray[14][19], Harray[15][19], Harray[16][19], Harray[17][19], Harray[18][19], Harray[19][19], Harray[20][19], Harray[21][19], Harray[22][19], Harray[23][19], Harray[24][19], Harray[25][19], Harray[26][19], Harray[27][19], Harray[28][19], Harray[29][19], Harray[30][19], Harray[31][19], Harray[32][19], Harray[33][19], Harray[34][19], Harray[35][19], Harray[36][19], Harray[37][19], Harray[38][19], Harray[39][19], Harray[40][19], Harray[41][19], Harray[42][19], Harray[43][19], Harray[44][19], Harray[45][19], Harray[46][19], Harray[47][19], Harray[48][19], Harray[49][19], Harray[50][19], Harray[51][19], Harray[52][19], Harray[53][19], Harray[54][19], Harray[55][19], Harray[56][19], Harray[57][19], Harray[58][19], Harray[59][19], Harray[60][19], Harray[61][19], Harray[62][19], Harray[63][19], Harray[64][19], Harray[65][19], Harray[66][19], Harray[67][19], Harray[68][19], Harray[69][19], Harray[70][19], Harray[71][19], Harray[72][19], Harray[73][19], Harray[74][19], Harray[75][19], Harray[76][19], Harray[77][19], Harray[78][19], Harray[79][19], Harray[80][19], Harray[81][19], Harray[82][19], Harray[83][19], Harray[84][19], Harray[85][19], Harray[86][19], Harray[87][19], Harray[88][19], Harray[89][19], Harray[90][19], Harray[91][19], Harray[92][19], Harray[93][19], Harray[94][19], Harray[95][19], Harray[96][19], Harray[97][19], Harray[98][19], Harray[99][19], Harray[100][19], Harray[101][19], Harray[102][19], Harray[103][19], Harray[104][19], Harray[105][19], Harray[106][19], Harray[107][19], Harray[108][19], Harray[109][19], Harray[110][19], Harray[111][19], Harray[112][19], Harray[113][19], Harray[114][19], Harray[115][19], Harray[116][19], Harray[117][19], Harray[118][19], Harray[119][19], Harray[120][19], Harray[121][19], Harray[122][19], Harray[123][19], Harray[124][19], Harray[125][19], Harray[126][19], Harray[127][19]};
assign h_col_20 = {Harray[0][20], Harray[1][20], Harray[2][20], Harray[3][20], Harray[4][20], Harray[5][20], Harray[6][20], Harray[7][20], Harray[8][20], Harray[9][20], Harray[10][20], Harray[11][20], Harray[12][20], Harray[13][20], Harray[14][20], Harray[15][20], Harray[16][20], Harray[17][20], Harray[18][20], Harray[19][20], Harray[20][20], Harray[21][20], Harray[22][20], Harray[23][20], Harray[24][20], Harray[25][20], Harray[26][20], Harray[27][20], Harray[28][20], Harray[29][20], Harray[30][20], Harray[31][20], Harray[32][20], Harray[33][20], Harray[34][20], Harray[35][20], Harray[36][20], Harray[37][20], Harray[38][20], Harray[39][20], Harray[40][20], Harray[41][20], Harray[42][20], Harray[43][20], Harray[44][20], Harray[45][20], Harray[46][20], Harray[47][20], Harray[48][20], Harray[49][20], Harray[50][20], Harray[51][20], Harray[52][20], Harray[53][20], Harray[54][20], Harray[55][20], Harray[56][20], Harray[57][20], Harray[58][20], Harray[59][20], Harray[60][20], Harray[61][20], Harray[62][20], Harray[63][20], Harray[64][20], Harray[65][20], Harray[66][20], Harray[67][20], Harray[68][20], Harray[69][20], Harray[70][20], Harray[71][20], Harray[72][20], Harray[73][20], Harray[74][20], Harray[75][20], Harray[76][20], Harray[77][20], Harray[78][20], Harray[79][20], Harray[80][20], Harray[81][20], Harray[82][20], Harray[83][20], Harray[84][20], Harray[85][20], Harray[86][20], Harray[87][20], Harray[88][20], Harray[89][20], Harray[90][20], Harray[91][20], Harray[92][20], Harray[93][20], Harray[94][20], Harray[95][20], Harray[96][20], Harray[97][20], Harray[98][20], Harray[99][20], Harray[100][20], Harray[101][20], Harray[102][20], Harray[103][20], Harray[104][20], Harray[105][20], Harray[106][20], Harray[107][20], Harray[108][20], Harray[109][20], Harray[110][20], Harray[111][20], Harray[112][20], Harray[113][20], Harray[114][20], Harray[115][20], Harray[116][20], Harray[117][20], Harray[118][20], Harray[119][20], Harray[120][20], Harray[121][20], Harray[122][20], Harray[123][20], Harray[124][20], Harray[125][20], Harray[126][20], Harray[127][20]};
assign h_col_21 = {Harray[0][21], Harray[1][21], Harray[2][21], Harray[3][21], Harray[4][21], Harray[5][21], Harray[6][21], Harray[7][21], Harray[8][21], Harray[9][21], Harray[10][21], Harray[11][21], Harray[12][21], Harray[13][21], Harray[14][21], Harray[15][21], Harray[16][21], Harray[17][21], Harray[18][21], Harray[19][21], Harray[20][21], Harray[21][21], Harray[22][21], Harray[23][21], Harray[24][21], Harray[25][21], Harray[26][21], Harray[27][21], Harray[28][21], Harray[29][21], Harray[30][21], Harray[31][21], Harray[32][21], Harray[33][21], Harray[34][21], Harray[35][21], Harray[36][21], Harray[37][21], Harray[38][21], Harray[39][21], Harray[40][21], Harray[41][21], Harray[42][21], Harray[43][21], Harray[44][21], Harray[45][21], Harray[46][21], Harray[47][21], Harray[48][21], Harray[49][21], Harray[50][21], Harray[51][21], Harray[52][21], Harray[53][21], Harray[54][21], Harray[55][21], Harray[56][21], Harray[57][21], Harray[58][21], Harray[59][21], Harray[60][21], Harray[61][21], Harray[62][21], Harray[63][21], Harray[64][21], Harray[65][21], Harray[66][21], Harray[67][21], Harray[68][21], Harray[69][21], Harray[70][21], Harray[71][21], Harray[72][21], Harray[73][21], Harray[74][21], Harray[75][21], Harray[76][21], Harray[77][21], Harray[78][21], Harray[79][21], Harray[80][21], Harray[81][21], Harray[82][21], Harray[83][21], Harray[84][21], Harray[85][21], Harray[86][21], Harray[87][21], Harray[88][21], Harray[89][21], Harray[90][21], Harray[91][21], Harray[92][21], Harray[93][21], Harray[94][21], Harray[95][21], Harray[96][21], Harray[97][21], Harray[98][21], Harray[99][21], Harray[100][21], Harray[101][21], Harray[102][21], Harray[103][21], Harray[104][21], Harray[105][21], Harray[106][21], Harray[107][21], Harray[108][21], Harray[109][21], Harray[110][21], Harray[111][21], Harray[112][21], Harray[113][21], Harray[114][21], Harray[115][21], Harray[116][21], Harray[117][21], Harray[118][21], Harray[119][21], Harray[120][21], Harray[121][21], Harray[122][21], Harray[123][21], Harray[124][21], Harray[125][21], Harray[126][21], Harray[127][21]};
assign h_col_22 = {Harray[0][22], Harray[1][22], Harray[2][22], Harray[3][22], Harray[4][22], Harray[5][22], Harray[6][22], Harray[7][22], Harray[8][22], Harray[9][22], Harray[10][22], Harray[11][22], Harray[12][22], Harray[13][22], Harray[14][22], Harray[15][22], Harray[16][22], Harray[17][22], Harray[18][22], Harray[19][22], Harray[20][22], Harray[21][22], Harray[22][22], Harray[23][22], Harray[24][22], Harray[25][22], Harray[26][22], Harray[27][22], Harray[28][22], Harray[29][22], Harray[30][22], Harray[31][22], Harray[32][22], Harray[33][22], Harray[34][22], Harray[35][22], Harray[36][22], Harray[37][22], Harray[38][22], Harray[39][22], Harray[40][22], Harray[41][22], Harray[42][22], Harray[43][22], Harray[44][22], Harray[45][22], Harray[46][22], Harray[47][22], Harray[48][22], Harray[49][22], Harray[50][22], Harray[51][22], Harray[52][22], Harray[53][22], Harray[54][22], Harray[55][22], Harray[56][22], Harray[57][22], Harray[58][22], Harray[59][22], Harray[60][22], Harray[61][22], Harray[62][22], Harray[63][22], Harray[64][22], Harray[65][22], Harray[66][22], Harray[67][22], Harray[68][22], Harray[69][22], Harray[70][22], Harray[71][22], Harray[72][22], Harray[73][22], Harray[74][22], Harray[75][22], Harray[76][22], Harray[77][22], Harray[78][22], Harray[79][22], Harray[80][22], Harray[81][22], Harray[82][22], Harray[83][22], Harray[84][22], Harray[85][22], Harray[86][22], Harray[87][22], Harray[88][22], Harray[89][22], Harray[90][22], Harray[91][22], Harray[92][22], Harray[93][22], Harray[94][22], Harray[95][22], Harray[96][22], Harray[97][22], Harray[98][22], Harray[99][22], Harray[100][22], Harray[101][22], Harray[102][22], Harray[103][22], Harray[104][22], Harray[105][22], Harray[106][22], Harray[107][22], Harray[108][22], Harray[109][22], Harray[110][22], Harray[111][22], Harray[112][22], Harray[113][22], Harray[114][22], Harray[115][22], Harray[116][22], Harray[117][22], Harray[118][22], Harray[119][22], Harray[120][22], Harray[121][22], Harray[122][22], Harray[123][22], Harray[124][22], Harray[125][22], Harray[126][22], Harray[127][22]};
assign h_col_23 = {Harray[0][23], Harray[1][23], Harray[2][23], Harray[3][23], Harray[4][23], Harray[5][23], Harray[6][23], Harray[7][23], Harray[8][23], Harray[9][23], Harray[10][23], Harray[11][23], Harray[12][23], Harray[13][23], Harray[14][23], Harray[15][23], Harray[16][23], Harray[17][23], Harray[18][23], Harray[19][23], Harray[20][23], Harray[21][23], Harray[22][23], Harray[23][23], Harray[24][23], Harray[25][23], Harray[26][23], Harray[27][23], Harray[28][23], Harray[29][23], Harray[30][23], Harray[31][23], Harray[32][23], Harray[33][23], Harray[34][23], Harray[35][23], Harray[36][23], Harray[37][23], Harray[38][23], Harray[39][23], Harray[40][23], Harray[41][23], Harray[42][23], Harray[43][23], Harray[44][23], Harray[45][23], Harray[46][23], Harray[47][23], Harray[48][23], Harray[49][23], Harray[50][23], Harray[51][23], Harray[52][23], Harray[53][23], Harray[54][23], Harray[55][23], Harray[56][23], Harray[57][23], Harray[58][23], Harray[59][23], Harray[60][23], Harray[61][23], Harray[62][23], Harray[63][23], Harray[64][23], Harray[65][23], Harray[66][23], Harray[67][23], Harray[68][23], Harray[69][23], Harray[70][23], Harray[71][23], Harray[72][23], Harray[73][23], Harray[74][23], Harray[75][23], Harray[76][23], Harray[77][23], Harray[78][23], Harray[79][23], Harray[80][23], Harray[81][23], Harray[82][23], Harray[83][23], Harray[84][23], Harray[85][23], Harray[86][23], Harray[87][23], Harray[88][23], Harray[89][23], Harray[90][23], Harray[91][23], Harray[92][23], Harray[93][23], Harray[94][23], Harray[95][23], Harray[96][23], Harray[97][23], Harray[98][23], Harray[99][23], Harray[100][23], Harray[101][23], Harray[102][23], Harray[103][23], Harray[104][23], Harray[105][23], Harray[106][23], Harray[107][23], Harray[108][23], Harray[109][23], Harray[110][23], Harray[111][23], Harray[112][23], Harray[113][23], Harray[114][23], Harray[115][23], Harray[116][23], Harray[117][23], Harray[118][23], Harray[119][23], Harray[120][23], Harray[121][23], Harray[122][23], Harray[123][23], Harray[124][23], Harray[125][23], Harray[126][23], Harray[127][23]};
assign h_col_24 = {Harray[0][24], Harray[1][24], Harray[2][24], Harray[3][24], Harray[4][24], Harray[5][24], Harray[6][24], Harray[7][24], Harray[8][24], Harray[9][24], Harray[10][24], Harray[11][24], Harray[12][24], Harray[13][24], Harray[14][24], Harray[15][24], Harray[16][24], Harray[17][24], Harray[18][24], Harray[19][24], Harray[20][24], Harray[21][24], Harray[22][24], Harray[23][24], Harray[24][24], Harray[25][24], Harray[26][24], Harray[27][24], Harray[28][24], Harray[29][24], Harray[30][24], Harray[31][24], Harray[32][24], Harray[33][24], Harray[34][24], Harray[35][24], Harray[36][24], Harray[37][24], Harray[38][24], Harray[39][24], Harray[40][24], Harray[41][24], Harray[42][24], Harray[43][24], Harray[44][24], Harray[45][24], Harray[46][24], Harray[47][24], Harray[48][24], Harray[49][24], Harray[50][24], Harray[51][24], Harray[52][24], Harray[53][24], Harray[54][24], Harray[55][24], Harray[56][24], Harray[57][24], Harray[58][24], Harray[59][24], Harray[60][24], Harray[61][24], Harray[62][24], Harray[63][24], Harray[64][24], Harray[65][24], Harray[66][24], Harray[67][24], Harray[68][24], Harray[69][24], Harray[70][24], Harray[71][24], Harray[72][24], Harray[73][24], Harray[74][24], Harray[75][24], Harray[76][24], Harray[77][24], Harray[78][24], Harray[79][24], Harray[80][24], Harray[81][24], Harray[82][24], Harray[83][24], Harray[84][24], Harray[85][24], Harray[86][24], Harray[87][24], Harray[88][24], Harray[89][24], Harray[90][24], Harray[91][24], Harray[92][24], Harray[93][24], Harray[94][24], Harray[95][24], Harray[96][24], Harray[97][24], Harray[98][24], Harray[99][24], Harray[100][24], Harray[101][24], Harray[102][24], Harray[103][24], Harray[104][24], Harray[105][24], Harray[106][24], Harray[107][24], Harray[108][24], Harray[109][24], Harray[110][24], Harray[111][24], Harray[112][24], Harray[113][24], Harray[114][24], Harray[115][24], Harray[116][24], Harray[117][24], Harray[118][24], Harray[119][24], Harray[120][24], Harray[121][24], Harray[122][24], Harray[123][24], Harray[124][24], Harray[125][24], Harray[126][24], Harray[127][24]};
assign h_col_25 = {Harray[0][25], Harray[1][25], Harray[2][25], Harray[3][25], Harray[4][25], Harray[5][25], Harray[6][25], Harray[7][25], Harray[8][25], Harray[9][25], Harray[10][25], Harray[11][25], Harray[12][25], Harray[13][25], Harray[14][25], Harray[15][25], Harray[16][25], Harray[17][25], Harray[18][25], Harray[19][25], Harray[20][25], Harray[21][25], Harray[22][25], Harray[23][25], Harray[24][25], Harray[25][25], Harray[26][25], Harray[27][25], Harray[28][25], Harray[29][25], Harray[30][25], Harray[31][25], Harray[32][25], Harray[33][25], Harray[34][25], Harray[35][25], Harray[36][25], Harray[37][25], Harray[38][25], Harray[39][25], Harray[40][25], Harray[41][25], Harray[42][25], Harray[43][25], Harray[44][25], Harray[45][25], Harray[46][25], Harray[47][25], Harray[48][25], Harray[49][25], Harray[50][25], Harray[51][25], Harray[52][25], Harray[53][25], Harray[54][25], Harray[55][25], Harray[56][25], Harray[57][25], Harray[58][25], Harray[59][25], Harray[60][25], Harray[61][25], Harray[62][25], Harray[63][25], Harray[64][25], Harray[65][25], Harray[66][25], Harray[67][25], Harray[68][25], Harray[69][25], Harray[70][25], Harray[71][25], Harray[72][25], Harray[73][25], Harray[74][25], Harray[75][25], Harray[76][25], Harray[77][25], Harray[78][25], Harray[79][25], Harray[80][25], Harray[81][25], Harray[82][25], Harray[83][25], Harray[84][25], Harray[85][25], Harray[86][25], Harray[87][25], Harray[88][25], Harray[89][25], Harray[90][25], Harray[91][25], Harray[92][25], Harray[93][25], Harray[94][25], Harray[95][25], Harray[96][25], Harray[97][25], Harray[98][25], Harray[99][25], Harray[100][25], Harray[101][25], Harray[102][25], Harray[103][25], Harray[104][25], Harray[105][25], Harray[106][25], Harray[107][25], Harray[108][25], Harray[109][25], Harray[110][25], Harray[111][25], Harray[112][25], Harray[113][25], Harray[114][25], Harray[115][25], Harray[116][25], Harray[117][25], Harray[118][25], Harray[119][25], Harray[120][25], Harray[121][25], Harray[122][25], Harray[123][25], Harray[124][25], Harray[125][25], Harray[126][25], Harray[127][25]};
assign h_col_26 = {Harray[0][26], Harray[1][26], Harray[2][26], Harray[3][26], Harray[4][26], Harray[5][26], Harray[6][26], Harray[7][26], Harray[8][26], Harray[9][26], Harray[10][26], Harray[11][26], Harray[12][26], Harray[13][26], Harray[14][26], Harray[15][26], Harray[16][26], Harray[17][26], Harray[18][26], Harray[19][26], Harray[20][26], Harray[21][26], Harray[22][26], Harray[23][26], Harray[24][26], Harray[25][26], Harray[26][26], Harray[27][26], Harray[28][26], Harray[29][26], Harray[30][26], Harray[31][26], Harray[32][26], Harray[33][26], Harray[34][26], Harray[35][26], Harray[36][26], Harray[37][26], Harray[38][26], Harray[39][26], Harray[40][26], Harray[41][26], Harray[42][26], Harray[43][26], Harray[44][26], Harray[45][26], Harray[46][26], Harray[47][26], Harray[48][26], Harray[49][26], Harray[50][26], Harray[51][26], Harray[52][26], Harray[53][26], Harray[54][26], Harray[55][26], Harray[56][26], Harray[57][26], Harray[58][26], Harray[59][26], Harray[60][26], Harray[61][26], Harray[62][26], Harray[63][26], Harray[64][26], Harray[65][26], Harray[66][26], Harray[67][26], Harray[68][26], Harray[69][26], Harray[70][26], Harray[71][26], Harray[72][26], Harray[73][26], Harray[74][26], Harray[75][26], Harray[76][26], Harray[77][26], Harray[78][26], Harray[79][26], Harray[80][26], Harray[81][26], Harray[82][26], Harray[83][26], Harray[84][26], Harray[85][26], Harray[86][26], Harray[87][26], Harray[88][26], Harray[89][26], Harray[90][26], Harray[91][26], Harray[92][26], Harray[93][26], Harray[94][26], Harray[95][26], Harray[96][26], Harray[97][26], Harray[98][26], Harray[99][26], Harray[100][26], Harray[101][26], Harray[102][26], Harray[103][26], Harray[104][26], Harray[105][26], Harray[106][26], Harray[107][26], Harray[108][26], Harray[109][26], Harray[110][26], Harray[111][26], Harray[112][26], Harray[113][26], Harray[114][26], Harray[115][26], Harray[116][26], Harray[117][26], Harray[118][26], Harray[119][26], Harray[120][26], Harray[121][26], Harray[122][26], Harray[123][26], Harray[124][26], Harray[125][26], Harray[126][26], Harray[127][26]};
assign h_col_27 = {Harray[0][27], Harray[1][27], Harray[2][27], Harray[3][27], Harray[4][27], Harray[5][27], Harray[6][27], Harray[7][27], Harray[8][27], Harray[9][27], Harray[10][27], Harray[11][27], Harray[12][27], Harray[13][27], Harray[14][27], Harray[15][27], Harray[16][27], Harray[17][27], Harray[18][27], Harray[19][27], Harray[20][27], Harray[21][27], Harray[22][27], Harray[23][27], Harray[24][27], Harray[25][27], Harray[26][27], Harray[27][27], Harray[28][27], Harray[29][27], Harray[30][27], Harray[31][27], Harray[32][27], Harray[33][27], Harray[34][27], Harray[35][27], Harray[36][27], Harray[37][27], Harray[38][27], Harray[39][27], Harray[40][27], Harray[41][27], Harray[42][27], Harray[43][27], Harray[44][27], Harray[45][27], Harray[46][27], Harray[47][27], Harray[48][27], Harray[49][27], Harray[50][27], Harray[51][27], Harray[52][27], Harray[53][27], Harray[54][27], Harray[55][27], Harray[56][27], Harray[57][27], Harray[58][27], Harray[59][27], Harray[60][27], Harray[61][27], Harray[62][27], Harray[63][27], Harray[64][27], Harray[65][27], Harray[66][27], Harray[67][27], Harray[68][27], Harray[69][27], Harray[70][27], Harray[71][27], Harray[72][27], Harray[73][27], Harray[74][27], Harray[75][27], Harray[76][27], Harray[77][27], Harray[78][27], Harray[79][27], Harray[80][27], Harray[81][27], Harray[82][27], Harray[83][27], Harray[84][27], Harray[85][27], Harray[86][27], Harray[87][27], Harray[88][27], Harray[89][27], Harray[90][27], Harray[91][27], Harray[92][27], Harray[93][27], Harray[94][27], Harray[95][27], Harray[96][27], Harray[97][27], Harray[98][27], Harray[99][27], Harray[100][27], Harray[101][27], Harray[102][27], Harray[103][27], Harray[104][27], Harray[105][27], Harray[106][27], Harray[107][27], Harray[108][27], Harray[109][27], Harray[110][27], Harray[111][27], Harray[112][27], Harray[113][27], Harray[114][27], Harray[115][27], Harray[116][27], Harray[117][27], Harray[118][27], Harray[119][27], Harray[120][27], Harray[121][27], Harray[122][27], Harray[123][27], Harray[124][27], Harray[125][27], Harray[126][27], Harray[127][27]};
assign h_col_28 = {Harray[0][28], Harray[1][28], Harray[2][28], Harray[3][28], Harray[4][28], Harray[5][28], Harray[6][28], Harray[7][28], Harray[8][28], Harray[9][28], Harray[10][28], Harray[11][28], Harray[12][28], Harray[13][28], Harray[14][28], Harray[15][28], Harray[16][28], Harray[17][28], Harray[18][28], Harray[19][28], Harray[20][28], Harray[21][28], Harray[22][28], Harray[23][28], Harray[24][28], Harray[25][28], Harray[26][28], Harray[27][28], Harray[28][28], Harray[29][28], Harray[30][28], Harray[31][28], Harray[32][28], Harray[33][28], Harray[34][28], Harray[35][28], Harray[36][28], Harray[37][28], Harray[38][28], Harray[39][28], Harray[40][28], Harray[41][28], Harray[42][28], Harray[43][28], Harray[44][28], Harray[45][28], Harray[46][28], Harray[47][28], Harray[48][28], Harray[49][28], Harray[50][28], Harray[51][28], Harray[52][28], Harray[53][28], Harray[54][28], Harray[55][28], Harray[56][28], Harray[57][28], Harray[58][28], Harray[59][28], Harray[60][28], Harray[61][28], Harray[62][28], Harray[63][28], Harray[64][28], Harray[65][28], Harray[66][28], Harray[67][28], Harray[68][28], Harray[69][28], Harray[70][28], Harray[71][28], Harray[72][28], Harray[73][28], Harray[74][28], Harray[75][28], Harray[76][28], Harray[77][28], Harray[78][28], Harray[79][28], Harray[80][28], Harray[81][28], Harray[82][28], Harray[83][28], Harray[84][28], Harray[85][28], Harray[86][28], Harray[87][28], Harray[88][28], Harray[89][28], Harray[90][28], Harray[91][28], Harray[92][28], Harray[93][28], Harray[94][28], Harray[95][28], Harray[96][28], Harray[97][28], Harray[98][28], Harray[99][28], Harray[100][28], Harray[101][28], Harray[102][28], Harray[103][28], Harray[104][28], Harray[105][28], Harray[106][28], Harray[107][28], Harray[108][28], Harray[109][28], Harray[110][28], Harray[111][28], Harray[112][28], Harray[113][28], Harray[114][28], Harray[115][28], Harray[116][28], Harray[117][28], Harray[118][28], Harray[119][28], Harray[120][28], Harray[121][28], Harray[122][28], Harray[123][28], Harray[124][28], Harray[125][28], Harray[126][28], Harray[127][28]};
assign h_col_29 = {Harray[0][29], Harray[1][29], Harray[2][29], Harray[3][29], Harray[4][29], Harray[5][29], Harray[6][29], Harray[7][29], Harray[8][29], Harray[9][29], Harray[10][29], Harray[11][29], Harray[12][29], Harray[13][29], Harray[14][29], Harray[15][29], Harray[16][29], Harray[17][29], Harray[18][29], Harray[19][29], Harray[20][29], Harray[21][29], Harray[22][29], Harray[23][29], Harray[24][29], Harray[25][29], Harray[26][29], Harray[27][29], Harray[28][29], Harray[29][29], Harray[30][29], Harray[31][29], Harray[32][29], Harray[33][29], Harray[34][29], Harray[35][29], Harray[36][29], Harray[37][29], Harray[38][29], Harray[39][29], Harray[40][29], Harray[41][29], Harray[42][29], Harray[43][29], Harray[44][29], Harray[45][29], Harray[46][29], Harray[47][29], Harray[48][29], Harray[49][29], Harray[50][29], Harray[51][29], Harray[52][29], Harray[53][29], Harray[54][29], Harray[55][29], Harray[56][29], Harray[57][29], Harray[58][29], Harray[59][29], Harray[60][29], Harray[61][29], Harray[62][29], Harray[63][29], Harray[64][29], Harray[65][29], Harray[66][29], Harray[67][29], Harray[68][29], Harray[69][29], Harray[70][29], Harray[71][29], Harray[72][29], Harray[73][29], Harray[74][29], Harray[75][29], Harray[76][29], Harray[77][29], Harray[78][29], Harray[79][29], Harray[80][29], Harray[81][29], Harray[82][29], Harray[83][29], Harray[84][29], Harray[85][29], Harray[86][29], Harray[87][29], Harray[88][29], Harray[89][29], Harray[90][29], Harray[91][29], Harray[92][29], Harray[93][29], Harray[94][29], Harray[95][29], Harray[96][29], Harray[97][29], Harray[98][29], Harray[99][29], Harray[100][29], Harray[101][29], Harray[102][29], Harray[103][29], Harray[104][29], Harray[105][29], Harray[106][29], Harray[107][29], Harray[108][29], Harray[109][29], Harray[110][29], Harray[111][29], Harray[112][29], Harray[113][29], Harray[114][29], Harray[115][29], Harray[116][29], Harray[117][29], Harray[118][29], Harray[119][29], Harray[120][29], Harray[121][29], Harray[122][29], Harray[123][29], Harray[124][29], Harray[125][29], Harray[126][29], Harray[127][29]};
assign h_col_30 = {Harray[0][30], Harray[1][30], Harray[2][30], Harray[3][30], Harray[4][30], Harray[5][30], Harray[6][30], Harray[7][30], Harray[8][30], Harray[9][30], Harray[10][30], Harray[11][30], Harray[12][30], Harray[13][30], Harray[14][30], Harray[15][30], Harray[16][30], Harray[17][30], Harray[18][30], Harray[19][30], Harray[20][30], Harray[21][30], Harray[22][30], Harray[23][30], Harray[24][30], Harray[25][30], Harray[26][30], Harray[27][30], Harray[28][30], Harray[29][30], Harray[30][30], Harray[31][30], Harray[32][30], Harray[33][30], Harray[34][30], Harray[35][30], Harray[36][30], Harray[37][30], Harray[38][30], Harray[39][30], Harray[40][30], Harray[41][30], Harray[42][30], Harray[43][30], Harray[44][30], Harray[45][30], Harray[46][30], Harray[47][30], Harray[48][30], Harray[49][30], Harray[50][30], Harray[51][30], Harray[52][30], Harray[53][30], Harray[54][30], Harray[55][30], Harray[56][30], Harray[57][30], Harray[58][30], Harray[59][30], Harray[60][30], Harray[61][30], Harray[62][30], Harray[63][30], Harray[64][30], Harray[65][30], Harray[66][30], Harray[67][30], Harray[68][30], Harray[69][30], Harray[70][30], Harray[71][30], Harray[72][30], Harray[73][30], Harray[74][30], Harray[75][30], Harray[76][30], Harray[77][30], Harray[78][30], Harray[79][30], Harray[80][30], Harray[81][30], Harray[82][30], Harray[83][30], Harray[84][30], Harray[85][30], Harray[86][30], Harray[87][30], Harray[88][30], Harray[89][30], Harray[90][30], Harray[91][30], Harray[92][30], Harray[93][30], Harray[94][30], Harray[95][30], Harray[96][30], Harray[97][30], Harray[98][30], Harray[99][30], Harray[100][30], Harray[101][30], Harray[102][30], Harray[103][30], Harray[104][30], Harray[105][30], Harray[106][30], Harray[107][30], Harray[108][30], Harray[109][30], Harray[110][30], Harray[111][30], Harray[112][30], Harray[113][30], Harray[114][30], Harray[115][30], Harray[116][30], Harray[117][30], Harray[118][30], Harray[119][30], Harray[120][30], Harray[121][30], Harray[122][30], Harray[123][30], Harray[124][30], Harray[125][30], Harray[126][30], Harray[127][30]};
assign h_col_31 = {Harray[0][31], Harray[1][31], Harray[2][31], Harray[3][31], Harray[4][31], Harray[5][31], Harray[6][31], Harray[7][31], Harray[8][31], Harray[9][31], Harray[10][31], Harray[11][31], Harray[12][31], Harray[13][31], Harray[14][31], Harray[15][31], Harray[16][31], Harray[17][31], Harray[18][31], Harray[19][31], Harray[20][31], Harray[21][31], Harray[22][31], Harray[23][31], Harray[24][31], Harray[25][31], Harray[26][31], Harray[27][31], Harray[28][31], Harray[29][31], Harray[30][31], Harray[31][31], Harray[32][31], Harray[33][31], Harray[34][31], Harray[35][31], Harray[36][31], Harray[37][31], Harray[38][31], Harray[39][31], Harray[40][31], Harray[41][31], Harray[42][31], Harray[43][31], Harray[44][31], Harray[45][31], Harray[46][31], Harray[47][31], Harray[48][31], Harray[49][31], Harray[50][31], Harray[51][31], Harray[52][31], Harray[53][31], Harray[54][31], Harray[55][31], Harray[56][31], Harray[57][31], Harray[58][31], Harray[59][31], Harray[60][31], Harray[61][31], Harray[62][31], Harray[63][31], Harray[64][31], Harray[65][31], Harray[66][31], Harray[67][31], Harray[68][31], Harray[69][31], Harray[70][31], Harray[71][31], Harray[72][31], Harray[73][31], Harray[74][31], Harray[75][31], Harray[76][31], Harray[77][31], Harray[78][31], Harray[79][31], Harray[80][31], Harray[81][31], Harray[82][31], Harray[83][31], Harray[84][31], Harray[85][31], Harray[86][31], Harray[87][31], Harray[88][31], Harray[89][31], Harray[90][31], Harray[91][31], Harray[92][31], Harray[93][31], Harray[94][31], Harray[95][31], Harray[96][31], Harray[97][31], Harray[98][31], Harray[99][31], Harray[100][31], Harray[101][31], Harray[102][31], Harray[103][31], Harray[104][31], Harray[105][31], Harray[106][31], Harray[107][31], Harray[108][31], Harray[109][31], Harray[110][31], Harray[111][31], Harray[112][31], Harray[113][31], Harray[114][31], Harray[115][31], Harray[116][31], Harray[117][31], Harray[118][31], Harray[119][31], Harray[120][31], Harray[121][31], Harray[122][31], Harray[123][31], Harray[124][31], Harray[125][31], Harray[126][31], Harray[127][31]};
assign h_col_32 = {Harray[0][32], Harray[1][32], Harray[2][32], Harray[3][32], Harray[4][32], Harray[5][32], Harray[6][32], Harray[7][32], Harray[8][32], Harray[9][32], Harray[10][32], Harray[11][32], Harray[12][32], Harray[13][32], Harray[14][32], Harray[15][32], Harray[16][32], Harray[17][32], Harray[18][32], Harray[19][32], Harray[20][32], Harray[21][32], Harray[22][32], Harray[23][32], Harray[24][32], Harray[25][32], Harray[26][32], Harray[27][32], Harray[28][32], Harray[29][32], Harray[30][32], Harray[31][32], Harray[32][32], Harray[33][32], Harray[34][32], Harray[35][32], Harray[36][32], Harray[37][32], Harray[38][32], Harray[39][32], Harray[40][32], Harray[41][32], Harray[42][32], Harray[43][32], Harray[44][32], Harray[45][32], Harray[46][32], Harray[47][32], Harray[48][32], Harray[49][32], Harray[50][32], Harray[51][32], Harray[52][32], Harray[53][32], Harray[54][32], Harray[55][32], Harray[56][32], Harray[57][32], Harray[58][32], Harray[59][32], Harray[60][32], Harray[61][32], Harray[62][32], Harray[63][32], Harray[64][32], Harray[65][32], Harray[66][32], Harray[67][32], Harray[68][32], Harray[69][32], Harray[70][32], Harray[71][32], Harray[72][32], Harray[73][32], Harray[74][32], Harray[75][32], Harray[76][32], Harray[77][32], Harray[78][32], Harray[79][32], Harray[80][32], Harray[81][32], Harray[82][32], Harray[83][32], Harray[84][32], Harray[85][32], Harray[86][32], Harray[87][32], Harray[88][32], Harray[89][32], Harray[90][32], Harray[91][32], Harray[92][32], Harray[93][32], Harray[94][32], Harray[95][32], Harray[96][32], Harray[97][32], Harray[98][32], Harray[99][32], Harray[100][32], Harray[101][32], Harray[102][32], Harray[103][32], Harray[104][32], Harray[105][32], Harray[106][32], Harray[107][32], Harray[108][32], Harray[109][32], Harray[110][32], Harray[111][32], Harray[112][32], Harray[113][32], Harray[114][32], Harray[115][32], Harray[116][32], Harray[117][32], Harray[118][32], Harray[119][32], Harray[120][32], Harray[121][32], Harray[122][32], Harray[123][32], Harray[124][32], Harray[125][32], Harray[126][32], Harray[127][32]};
assign h_col_33 = {Harray[0][33], Harray[1][33], Harray[2][33], Harray[3][33], Harray[4][33], Harray[5][33], Harray[6][33], Harray[7][33], Harray[8][33], Harray[9][33], Harray[10][33], Harray[11][33], Harray[12][33], Harray[13][33], Harray[14][33], Harray[15][33], Harray[16][33], Harray[17][33], Harray[18][33], Harray[19][33], Harray[20][33], Harray[21][33], Harray[22][33], Harray[23][33], Harray[24][33], Harray[25][33], Harray[26][33], Harray[27][33], Harray[28][33], Harray[29][33], Harray[30][33], Harray[31][33], Harray[32][33], Harray[33][33], Harray[34][33], Harray[35][33], Harray[36][33], Harray[37][33], Harray[38][33], Harray[39][33], Harray[40][33], Harray[41][33], Harray[42][33], Harray[43][33], Harray[44][33], Harray[45][33], Harray[46][33], Harray[47][33], Harray[48][33], Harray[49][33], Harray[50][33], Harray[51][33], Harray[52][33], Harray[53][33], Harray[54][33], Harray[55][33], Harray[56][33], Harray[57][33], Harray[58][33], Harray[59][33], Harray[60][33], Harray[61][33], Harray[62][33], Harray[63][33], Harray[64][33], Harray[65][33], Harray[66][33], Harray[67][33], Harray[68][33], Harray[69][33], Harray[70][33], Harray[71][33], Harray[72][33], Harray[73][33], Harray[74][33], Harray[75][33], Harray[76][33], Harray[77][33], Harray[78][33], Harray[79][33], Harray[80][33], Harray[81][33], Harray[82][33], Harray[83][33], Harray[84][33], Harray[85][33], Harray[86][33], Harray[87][33], Harray[88][33], Harray[89][33], Harray[90][33], Harray[91][33], Harray[92][33], Harray[93][33], Harray[94][33], Harray[95][33], Harray[96][33], Harray[97][33], Harray[98][33], Harray[99][33], Harray[100][33], Harray[101][33], Harray[102][33], Harray[103][33], Harray[104][33], Harray[105][33], Harray[106][33], Harray[107][33], Harray[108][33], Harray[109][33], Harray[110][33], Harray[111][33], Harray[112][33], Harray[113][33], Harray[114][33], Harray[115][33], Harray[116][33], Harray[117][33], Harray[118][33], Harray[119][33], Harray[120][33], Harray[121][33], Harray[122][33], Harray[123][33], Harray[124][33], Harray[125][33], Harray[126][33], Harray[127][33]};
assign h_col_34 = {Harray[0][34], Harray[1][34], Harray[2][34], Harray[3][34], Harray[4][34], Harray[5][34], Harray[6][34], Harray[7][34], Harray[8][34], Harray[9][34], Harray[10][34], Harray[11][34], Harray[12][34], Harray[13][34], Harray[14][34], Harray[15][34], Harray[16][34], Harray[17][34], Harray[18][34], Harray[19][34], Harray[20][34], Harray[21][34], Harray[22][34], Harray[23][34], Harray[24][34], Harray[25][34], Harray[26][34], Harray[27][34], Harray[28][34], Harray[29][34], Harray[30][34], Harray[31][34], Harray[32][34], Harray[33][34], Harray[34][34], Harray[35][34], Harray[36][34], Harray[37][34], Harray[38][34], Harray[39][34], Harray[40][34], Harray[41][34], Harray[42][34], Harray[43][34], Harray[44][34], Harray[45][34], Harray[46][34], Harray[47][34], Harray[48][34], Harray[49][34], Harray[50][34], Harray[51][34], Harray[52][34], Harray[53][34], Harray[54][34], Harray[55][34], Harray[56][34], Harray[57][34], Harray[58][34], Harray[59][34], Harray[60][34], Harray[61][34], Harray[62][34], Harray[63][34], Harray[64][34], Harray[65][34], Harray[66][34], Harray[67][34], Harray[68][34], Harray[69][34], Harray[70][34], Harray[71][34], Harray[72][34], Harray[73][34], Harray[74][34], Harray[75][34], Harray[76][34], Harray[77][34], Harray[78][34], Harray[79][34], Harray[80][34], Harray[81][34], Harray[82][34], Harray[83][34], Harray[84][34], Harray[85][34], Harray[86][34], Harray[87][34], Harray[88][34], Harray[89][34], Harray[90][34], Harray[91][34], Harray[92][34], Harray[93][34], Harray[94][34], Harray[95][34], Harray[96][34], Harray[97][34], Harray[98][34], Harray[99][34], Harray[100][34], Harray[101][34], Harray[102][34], Harray[103][34], Harray[104][34], Harray[105][34], Harray[106][34], Harray[107][34], Harray[108][34], Harray[109][34], Harray[110][34], Harray[111][34], Harray[112][34], Harray[113][34], Harray[114][34], Harray[115][34], Harray[116][34], Harray[117][34], Harray[118][34], Harray[119][34], Harray[120][34], Harray[121][34], Harray[122][34], Harray[123][34], Harray[124][34], Harray[125][34], Harray[126][34], Harray[127][34]};
assign h_col_35 = {Harray[0][35], Harray[1][35], Harray[2][35], Harray[3][35], Harray[4][35], Harray[5][35], Harray[6][35], Harray[7][35], Harray[8][35], Harray[9][35], Harray[10][35], Harray[11][35], Harray[12][35], Harray[13][35], Harray[14][35], Harray[15][35], Harray[16][35], Harray[17][35], Harray[18][35], Harray[19][35], Harray[20][35], Harray[21][35], Harray[22][35], Harray[23][35], Harray[24][35], Harray[25][35], Harray[26][35], Harray[27][35], Harray[28][35], Harray[29][35], Harray[30][35], Harray[31][35], Harray[32][35], Harray[33][35], Harray[34][35], Harray[35][35], Harray[36][35], Harray[37][35], Harray[38][35], Harray[39][35], Harray[40][35], Harray[41][35], Harray[42][35], Harray[43][35], Harray[44][35], Harray[45][35], Harray[46][35], Harray[47][35], Harray[48][35], Harray[49][35], Harray[50][35], Harray[51][35], Harray[52][35], Harray[53][35], Harray[54][35], Harray[55][35], Harray[56][35], Harray[57][35], Harray[58][35], Harray[59][35], Harray[60][35], Harray[61][35], Harray[62][35], Harray[63][35], Harray[64][35], Harray[65][35], Harray[66][35], Harray[67][35], Harray[68][35], Harray[69][35], Harray[70][35], Harray[71][35], Harray[72][35], Harray[73][35], Harray[74][35], Harray[75][35], Harray[76][35], Harray[77][35], Harray[78][35], Harray[79][35], Harray[80][35], Harray[81][35], Harray[82][35], Harray[83][35], Harray[84][35], Harray[85][35], Harray[86][35], Harray[87][35], Harray[88][35], Harray[89][35], Harray[90][35], Harray[91][35], Harray[92][35], Harray[93][35], Harray[94][35], Harray[95][35], Harray[96][35], Harray[97][35], Harray[98][35], Harray[99][35], Harray[100][35], Harray[101][35], Harray[102][35], Harray[103][35], Harray[104][35], Harray[105][35], Harray[106][35], Harray[107][35], Harray[108][35], Harray[109][35], Harray[110][35], Harray[111][35], Harray[112][35], Harray[113][35], Harray[114][35], Harray[115][35], Harray[116][35], Harray[117][35], Harray[118][35], Harray[119][35], Harray[120][35], Harray[121][35], Harray[122][35], Harray[123][35], Harray[124][35], Harray[125][35], Harray[126][35], Harray[127][35]};
assign h_col_36 = {Harray[0][36], Harray[1][36], Harray[2][36], Harray[3][36], Harray[4][36], Harray[5][36], Harray[6][36], Harray[7][36], Harray[8][36], Harray[9][36], Harray[10][36], Harray[11][36], Harray[12][36], Harray[13][36], Harray[14][36], Harray[15][36], Harray[16][36], Harray[17][36], Harray[18][36], Harray[19][36], Harray[20][36], Harray[21][36], Harray[22][36], Harray[23][36], Harray[24][36], Harray[25][36], Harray[26][36], Harray[27][36], Harray[28][36], Harray[29][36], Harray[30][36], Harray[31][36], Harray[32][36], Harray[33][36], Harray[34][36], Harray[35][36], Harray[36][36], Harray[37][36], Harray[38][36], Harray[39][36], Harray[40][36], Harray[41][36], Harray[42][36], Harray[43][36], Harray[44][36], Harray[45][36], Harray[46][36], Harray[47][36], Harray[48][36], Harray[49][36], Harray[50][36], Harray[51][36], Harray[52][36], Harray[53][36], Harray[54][36], Harray[55][36], Harray[56][36], Harray[57][36], Harray[58][36], Harray[59][36], Harray[60][36], Harray[61][36], Harray[62][36], Harray[63][36], Harray[64][36], Harray[65][36], Harray[66][36], Harray[67][36], Harray[68][36], Harray[69][36], Harray[70][36], Harray[71][36], Harray[72][36], Harray[73][36], Harray[74][36], Harray[75][36], Harray[76][36], Harray[77][36], Harray[78][36], Harray[79][36], Harray[80][36], Harray[81][36], Harray[82][36], Harray[83][36], Harray[84][36], Harray[85][36], Harray[86][36], Harray[87][36], Harray[88][36], Harray[89][36], Harray[90][36], Harray[91][36], Harray[92][36], Harray[93][36], Harray[94][36], Harray[95][36], Harray[96][36], Harray[97][36], Harray[98][36], Harray[99][36], Harray[100][36], Harray[101][36], Harray[102][36], Harray[103][36], Harray[104][36], Harray[105][36], Harray[106][36], Harray[107][36], Harray[108][36], Harray[109][36], Harray[110][36], Harray[111][36], Harray[112][36], Harray[113][36], Harray[114][36], Harray[115][36], Harray[116][36], Harray[117][36], Harray[118][36], Harray[119][36], Harray[120][36], Harray[121][36], Harray[122][36], Harray[123][36], Harray[124][36], Harray[125][36], Harray[126][36], Harray[127][36]};
assign h_col_37 = {Harray[0][37], Harray[1][37], Harray[2][37], Harray[3][37], Harray[4][37], Harray[5][37], Harray[6][37], Harray[7][37], Harray[8][37], Harray[9][37], Harray[10][37], Harray[11][37], Harray[12][37], Harray[13][37], Harray[14][37], Harray[15][37], Harray[16][37], Harray[17][37], Harray[18][37], Harray[19][37], Harray[20][37], Harray[21][37], Harray[22][37], Harray[23][37], Harray[24][37], Harray[25][37], Harray[26][37], Harray[27][37], Harray[28][37], Harray[29][37], Harray[30][37], Harray[31][37], Harray[32][37], Harray[33][37], Harray[34][37], Harray[35][37], Harray[36][37], Harray[37][37], Harray[38][37], Harray[39][37], Harray[40][37], Harray[41][37], Harray[42][37], Harray[43][37], Harray[44][37], Harray[45][37], Harray[46][37], Harray[47][37], Harray[48][37], Harray[49][37], Harray[50][37], Harray[51][37], Harray[52][37], Harray[53][37], Harray[54][37], Harray[55][37], Harray[56][37], Harray[57][37], Harray[58][37], Harray[59][37], Harray[60][37], Harray[61][37], Harray[62][37], Harray[63][37], Harray[64][37], Harray[65][37], Harray[66][37], Harray[67][37], Harray[68][37], Harray[69][37], Harray[70][37], Harray[71][37], Harray[72][37], Harray[73][37], Harray[74][37], Harray[75][37], Harray[76][37], Harray[77][37], Harray[78][37], Harray[79][37], Harray[80][37], Harray[81][37], Harray[82][37], Harray[83][37], Harray[84][37], Harray[85][37], Harray[86][37], Harray[87][37], Harray[88][37], Harray[89][37], Harray[90][37], Harray[91][37], Harray[92][37], Harray[93][37], Harray[94][37], Harray[95][37], Harray[96][37], Harray[97][37], Harray[98][37], Harray[99][37], Harray[100][37], Harray[101][37], Harray[102][37], Harray[103][37], Harray[104][37], Harray[105][37], Harray[106][37], Harray[107][37], Harray[108][37], Harray[109][37], Harray[110][37], Harray[111][37], Harray[112][37], Harray[113][37], Harray[114][37], Harray[115][37], Harray[116][37], Harray[117][37], Harray[118][37], Harray[119][37], Harray[120][37], Harray[121][37], Harray[122][37], Harray[123][37], Harray[124][37], Harray[125][37], Harray[126][37], Harray[127][37]};
assign h_col_38 = {Harray[0][38], Harray[1][38], Harray[2][38], Harray[3][38], Harray[4][38], Harray[5][38], Harray[6][38], Harray[7][38], Harray[8][38], Harray[9][38], Harray[10][38], Harray[11][38], Harray[12][38], Harray[13][38], Harray[14][38], Harray[15][38], Harray[16][38], Harray[17][38], Harray[18][38], Harray[19][38], Harray[20][38], Harray[21][38], Harray[22][38], Harray[23][38], Harray[24][38], Harray[25][38], Harray[26][38], Harray[27][38], Harray[28][38], Harray[29][38], Harray[30][38], Harray[31][38], Harray[32][38], Harray[33][38], Harray[34][38], Harray[35][38], Harray[36][38], Harray[37][38], Harray[38][38], Harray[39][38], Harray[40][38], Harray[41][38], Harray[42][38], Harray[43][38], Harray[44][38], Harray[45][38], Harray[46][38], Harray[47][38], Harray[48][38], Harray[49][38], Harray[50][38], Harray[51][38], Harray[52][38], Harray[53][38], Harray[54][38], Harray[55][38], Harray[56][38], Harray[57][38], Harray[58][38], Harray[59][38], Harray[60][38], Harray[61][38], Harray[62][38], Harray[63][38], Harray[64][38], Harray[65][38], Harray[66][38], Harray[67][38], Harray[68][38], Harray[69][38], Harray[70][38], Harray[71][38], Harray[72][38], Harray[73][38], Harray[74][38], Harray[75][38], Harray[76][38], Harray[77][38], Harray[78][38], Harray[79][38], Harray[80][38], Harray[81][38], Harray[82][38], Harray[83][38], Harray[84][38], Harray[85][38], Harray[86][38], Harray[87][38], Harray[88][38], Harray[89][38], Harray[90][38], Harray[91][38], Harray[92][38], Harray[93][38], Harray[94][38], Harray[95][38], Harray[96][38], Harray[97][38], Harray[98][38], Harray[99][38], Harray[100][38], Harray[101][38], Harray[102][38], Harray[103][38], Harray[104][38], Harray[105][38], Harray[106][38], Harray[107][38], Harray[108][38], Harray[109][38], Harray[110][38], Harray[111][38], Harray[112][38], Harray[113][38], Harray[114][38], Harray[115][38], Harray[116][38], Harray[117][38], Harray[118][38], Harray[119][38], Harray[120][38], Harray[121][38], Harray[122][38], Harray[123][38], Harray[124][38], Harray[125][38], Harray[126][38], Harray[127][38]};
assign h_col_39 = {Harray[0][39], Harray[1][39], Harray[2][39], Harray[3][39], Harray[4][39], Harray[5][39], Harray[6][39], Harray[7][39], Harray[8][39], Harray[9][39], Harray[10][39], Harray[11][39], Harray[12][39], Harray[13][39], Harray[14][39], Harray[15][39], Harray[16][39], Harray[17][39], Harray[18][39], Harray[19][39], Harray[20][39], Harray[21][39], Harray[22][39], Harray[23][39], Harray[24][39], Harray[25][39], Harray[26][39], Harray[27][39], Harray[28][39], Harray[29][39], Harray[30][39], Harray[31][39], Harray[32][39], Harray[33][39], Harray[34][39], Harray[35][39], Harray[36][39], Harray[37][39], Harray[38][39], Harray[39][39], Harray[40][39], Harray[41][39], Harray[42][39], Harray[43][39], Harray[44][39], Harray[45][39], Harray[46][39], Harray[47][39], Harray[48][39], Harray[49][39], Harray[50][39], Harray[51][39], Harray[52][39], Harray[53][39], Harray[54][39], Harray[55][39], Harray[56][39], Harray[57][39], Harray[58][39], Harray[59][39], Harray[60][39], Harray[61][39], Harray[62][39], Harray[63][39], Harray[64][39], Harray[65][39], Harray[66][39], Harray[67][39], Harray[68][39], Harray[69][39], Harray[70][39], Harray[71][39], Harray[72][39], Harray[73][39], Harray[74][39], Harray[75][39], Harray[76][39], Harray[77][39], Harray[78][39], Harray[79][39], Harray[80][39], Harray[81][39], Harray[82][39], Harray[83][39], Harray[84][39], Harray[85][39], Harray[86][39], Harray[87][39], Harray[88][39], Harray[89][39], Harray[90][39], Harray[91][39], Harray[92][39], Harray[93][39], Harray[94][39], Harray[95][39], Harray[96][39], Harray[97][39], Harray[98][39], Harray[99][39], Harray[100][39], Harray[101][39], Harray[102][39], Harray[103][39], Harray[104][39], Harray[105][39], Harray[106][39], Harray[107][39], Harray[108][39], Harray[109][39], Harray[110][39], Harray[111][39], Harray[112][39], Harray[113][39], Harray[114][39], Harray[115][39], Harray[116][39], Harray[117][39], Harray[118][39], Harray[119][39], Harray[120][39], Harray[121][39], Harray[122][39], Harray[123][39], Harray[124][39], Harray[125][39], Harray[126][39], Harray[127][39]};
assign h_col_40 = {Harray[0][40], Harray[1][40], Harray[2][40], Harray[3][40], Harray[4][40], Harray[5][40], Harray[6][40], Harray[7][40], Harray[8][40], Harray[9][40], Harray[10][40], Harray[11][40], Harray[12][40], Harray[13][40], Harray[14][40], Harray[15][40], Harray[16][40], Harray[17][40], Harray[18][40], Harray[19][40], Harray[20][40], Harray[21][40], Harray[22][40], Harray[23][40], Harray[24][40], Harray[25][40], Harray[26][40], Harray[27][40], Harray[28][40], Harray[29][40], Harray[30][40], Harray[31][40], Harray[32][40], Harray[33][40], Harray[34][40], Harray[35][40], Harray[36][40], Harray[37][40], Harray[38][40], Harray[39][40], Harray[40][40], Harray[41][40], Harray[42][40], Harray[43][40], Harray[44][40], Harray[45][40], Harray[46][40], Harray[47][40], Harray[48][40], Harray[49][40], Harray[50][40], Harray[51][40], Harray[52][40], Harray[53][40], Harray[54][40], Harray[55][40], Harray[56][40], Harray[57][40], Harray[58][40], Harray[59][40], Harray[60][40], Harray[61][40], Harray[62][40], Harray[63][40], Harray[64][40], Harray[65][40], Harray[66][40], Harray[67][40], Harray[68][40], Harray[69][40], Harray[70][40], Harray[71][40], Harray[72][40], Harray[73][40], Harray[74][40], Harray[75][40], Harray[76][40], Harray[77][40], Harray[78][40], Harray[79][40], Harray[80][40], Harray[81][40], Harray[82][40], Harray[83][40], Harray[84][40], Harray[85][40], Harray[86][40], Harray[87][40], Harray[88][40], Harray[89][40], Harray[90][40], Harray[91][40], Harray[92][40], Harray[93][40], Harray[94][40], Harray[95][40], Harray[96][40], Harray[97][40], Harray[98][40], Harray[99][40], Harray[100][40], Harray[101][40], Harray[102][40], Harray[103][40], Harray[104][40], Harray[105][40], Harray[106][40], Harray[107][40], Harray[108][40], Harray[109][40], Harray[110][40], Harray[111][40], Harray[112][40], Harray[113][40], Harray[114][40], Harray[115][40], Harray[116][40], Harray[117][40], Harray[118][40], Harray[119][40], Harray[120][40], Harray[121][40], Harray[122][40], Harray[123][40], Harray[124][40], Harray[125][40], Harray[126][40], Harray[127][40]};
assign h_col_41 = {Harray[0][41], Harray[1][41], Harray[2][41], Harray[3][41], Harray[4][41], Harray[5][41], Harray[6][41], Harray[7][41], Harray[8][41], Harray[9][41], Harray[10][41], Harray[11][41], Harray[12][41], Harray[13][41], Harray[14][41], Harray[15][41], Harray[16][41], Harray[17][41], Harray[18][41], Harray[19][41], Harray[20][41], Harray[21][41], Harray[22][41], Harray[23][41], Harray[24][41], Harray[25][41], Harray[26][41], Harray[27][41], Harray[28][41], Harray[29][41], Harray[30][41], Harray[31][41], Harray[32][41], Harray[33][41], Harray[34][41], Harray[35][41], Harray[36][41], Harray[37][41], Harray[38][41], Harray[39][41], Harray[40][41], Harray[41][41], Harray[42][41], Harray[43][41], Harray[44][41], Harray[45][41], Harray[46][41], Harray[47][41], Harray[48][41], Harray[49][41], Harray[50][41], Harray[51][41], Harray[52][41], Harray[53][41], Harray[54][41], Harray[55][41], Harray[56][41], Harray[57][41], Harray[58][41], Harray[59][41], Harray[60][41], Harray[61][41], Harray[62][41], Harray[63][41], Harray[64][41], Harray[65][41], Harray[66][41], Harray[67][41], Harray[68][41], Harray[69][41], Harray[70][41], Harray[71][41], Harray[72][41], Harray[73][41], Harray[74][41], Harray[75][41], Harray[76][41], Harray[77][41], Harray[78][41], Harray[79][41], Harray[80][41], Harray[81][41], Harray[82][41], Harray[83][41], Harray[84][41], Harray[85][41], Harray[86][41], Harray[87][41], Harray[88][41], Harray[89][41], Harray[90][41], Harray[91][41], Harray[92][41], Harray[93][41], Harray[94][41], Harray[95][41], Harray[96][41], Harray[97][41], Harray[98][41], Harray[99][41], Harray[100][41], Harray[101][41], Harray[102][41], Harray[103][41], Harray[104][41], Harray[105][41], Harray[106][41], Harray[107][41], Harray[108][41], Harray[109][41], Harray[110][41], Harray[111][41], Harray[112][41], Harray[113][41], Harray[114][41], Harray[115][41], Harray[116][41], Harray[117][41], Harray[118][41], Harray[119][41], Harray[120][41], Harray[121][41], Harray[122][41], Harray[123][41], Harray[124][41], Harray[125][41], Harray[126][41], Harray[127][41]};
assign h_col_42 = {Harray[0][42], Harray[1][42], Harray[2][42], Harray[3][42], Harray[4][42], Harray[5][42], Harray[6][42], Harray[7][42], Harray[8][42], Harray[9][42], Harray[10][42], Harray[11][42], Harray[12][42], Harray[13][42], Harray[14][42], Harray[15][42], Harray[16][42], Harray[17][42], Harray[18][42], Harray[19][42], Harray[20][42], Harray[21][42], Harray[22][42], Harray[23][42], Harray[24][42], Harray[25][42], Harray[26][42], Harray[27][42], Harray[28][42], Harray[29][42], Harray[30][42], Harray[31][42], Harray[32][42], Harray[33][42], Harray[34][42], Harray[35][42], Harray[36][42], Harray[37][42], Harray[38][42], Harray[39][42], Harray[40][42], Harray[41][42], Harray[42][42], Harray[43][42], Harray[44][42], Harray[45][42], Harray[46][42], Harray[47][42], Harray[48][42], Harray[49][42], Harray[50][42], Harray[51][42], Harray[52][42], Harray[53][42], Harray[54][42], Harray[55][42], Harray[56][42], Harray[57][42], Harray[58][42], Harray[59][42], Harray[60][42], Harray[61][42], Harray[62][42], Harray[63][42], Harray[64][42], Harray[65][42], Harray[66][42], Harray[67][42], Harray[68][42], Harray[69][42], Harray[70][42], Harray[71][42], Harray[72][42], Harray[73][42], Harray[74][42], Harray[75][42], Harray[76][42], Harray[77][42], Harray[78][42], Harray[79][42], Harray[80][42], Harray[81][42], Harray[82][42], Harray[83][42], Harray[84][42], Harray[85][42], Harray[86][42], Harray[87][42], Harray[88][42], Harray[89][42], Harray[90][42], Harray[91][42], Harray[92][42], Harray[93][42], Harray[94][42], Harray[95][42], Harray[96][42], Harray[97][42], Harray[98][42], Harray[99][42], Harray[100][42], Harray[101][42], Harray[102][42], Harray[103][42], Harray[104][42], Harray[105][42], Harray[106][42], Harray[107][42], Harray[108][42], Harray[109][42], Harray[110][42], Harray[111][42], Harray[112][42], Harray[113][42], Harray[114][42], Harray[115][42], Harray[116][42], Harray[117][42], Harray[118][42], Harray[119][42], Harray[120][42], Harray[121][42], Harray[122][42], Harray[123][42], Harray[124][42], Harray[125][42], Harray[126][42], Harray[127][42]};
assign h_col_43 = {Harray[0][43], Harray[1][43], Harray[2][43], Harray[3][43], Harray[4][43], Harray[5][43], Harray[6][43], Harray[7][43], Harray[8][43], Harray[9][43], Harray[10][43], Harray[11][43], Harray[12][43], Harray[13][43], Harray[14][43], Harray[15][43], Harray[16][43], Harray[17][43], Harray[18][43], Harray[19][43], Harray[20][43], Harray[21][43], Harray[22][43], Harray[23][43], Harray[24][43], Harray[25][43], Harray[26][43], Harray[27][43], Harray[28][43], Harray[29][43], Harray[30][43], Harray[31][43], Harray[32][43], Harray[33][43], Harray[34][43], Harray[35][43], Harray[36][43], Harray[37][43], Harray[38][43], Harray[39][43], Harray[40][43], Harray[41][43], Harray[42][43], Harray[43][43], Harray[44][43], Harray[45][43], Harray[46][43], Harray[47][43], Harray[48][43], Harray[49][43], Harray[50][43], Harray[51][43], Harray[52][43], Harray[53][43], Harray[54][43], Harray[55][43], Harray[56][43], Harray[57][43], Harray[58][43], Harray[59][43], Harray[60][43], Harray[61][43], Harray[62][43], Harray[63][43], Harray[64][43], Harray[65][43], Harray[66][43], Harray[67][43], Harray[68][43], Harray[69][43], Harray[70][43], Harray[71][43], Harray[72][43], Harray[73][43], Harray[74][43], Harray[75][43], Harray[76][43], Harray[77][43], Harray[78][43], Harray[79][43], Harray[80][43], Harray[81][43], Harray[82][43], Harray[83][43], Harray[84][43], Harray[85][43], Harray[86][43], Harray[87][43], Harray[88][43], Harray[89][43], Harray[90][43], Harray[91][43], Harray[92][43], Harray[93][43], Harray[94][43], Harray[95][43], Harray[96][43], Harray[97][43], Harray[98][43], Harray[99][43], Harray[100][43], Harray[101][43], Harray[102][43], Harray[103][43], Harray[104][43], Harray[105][43], Harray[106][43], Harray[107][43], Harray[108][43], Harray[109][43], Harray[110][43], Harray[111][43], Harray[112][43], Harray[113][43], Harray[114][43], Harray[115][43], Harray[116][43], Harray[117][43], Harray[118][43], Harray[119][43], Harray[120][43], Harray[121][43], Harray[122][43], Harray[123][43], Harray[124][43], Harray[125][43], Harray[126][43], Harray[127][43]};
assign h_col_44 = {Harray[0][44], Harray[1][44], Harray[2][44], Harray[3][44], Harray[4][44], Harray[5][44], Harray[6][44], Harray[7][44], Harray[8][44], Harray[9][44], Harray[10][44], Harray[11][44], Harray[12][44], Harray[13][44], Harray[14][44], Harray[15][44], Harray[16][44], Harray[17][44], Harray[18][44], Harray[19][44], Harray[20][44], Harray[21][44], Harray[22][44], Harray[23][44], Harray[24][44], Harray[25][44], Harray[26][44], Harray[27][44], Harray[28][44], Harray[29][44], Harray[30][44], Harray[31][44], Harray[32][44], Harray[33][44], Harray[34][44], Harray[35][44], Harray[36][44], Harray[37][44], Harray[38][44], Harray[39][44], Harray[40][44], Harray[41][44], Harray[42][44], Harray[43][44], Harray[44][44], Harray[45][44], Harray[46][44], Harray[47][44], Harray[48][44], Harray[49][44], Harray[50][44], Harray[51][44], Harray[52][44], Harray[53][44], Harray[54][44], Harray[55][44], Harray[56][44], Harray[57][44], Harray[58][44], Harray[59][44], Harray[60][44], Harray[61][44], Harray[62][44], Harray[63][44], Harray[64][44], Harray[65][44], Harray[66][44], Harray[67][44], Harray[68][44], Harray[69][44], Harray[70][44], Harray[71][44], Harray[72][44], Harray[73][44], Harray[74][44], Harray[75][44], Harray[76][44], Harray[77][44], Harray[78][44], Harray[79][44], Harray[80][44], Harray[81][44], Harray[82][44], Harray[83][44], Harray[84][44], Harray[85][44], Harray[86][44], Harray[87][44], Harray[88][44], Harray[89][44], Harray[90][44], Harray[91][44], Harray[92][44], Harray[93][44], Harray[94][44], Harray[95][44], Harray[96][44], Harray[97][44], Harray[98][44], Harray[99][44], Harray[100][44], Harray[101][44], Harray[102][44], Harray[103][44], Harray[104][44], Harray[105][44], Harray[106][44], Harray[107][44], Harray[108][44], Harray[109][44], Harray[110][44], Harray[111][44], Harray[112][44], Harray[113][44], Harray[114][44], Harray[115][44], Harray[116][44], Harray[117][44], Harray[118][44], Harray[119][44], Harray[120][44], Harray[121][44], Harray[122][44], Harray[123][44], Harray[124][44], Harray[125][44], Harray[126][44], Harray[127][44]};
assign h_col_45 = {Harray[0][45], Harray[1][45], Harray[2][45], Harray[3][45], Harray[4][45], Harray[5][45], Harray[6][45], Harray[7][45], Harray[8][45], Harray[9][45], Harray[10][45], Harray[11][45], Harray[12][45], Harray[13][45], Harray[14][45], Harray[15][45], Harray[16][45], Harray[17][45], Harray[18][45], Harray[19][45], Harray[20][45], Harray[21][45], Harray[22][45], Harray[23][45], Harray[24][45], Harray[25][45], Harray[26][45], Harray[27][45], Harray[28][45], Harray[29][45], Harray[30][45], Harray[31][45], Harray[32][45], Harray[33][45], Harray[34][45], Harray[35][45], Harray[36][45], Harray[37][45], Harray[38][45], Harray[39][45], Harray[40][45], Harray[41][45], Harray[42][45], Harray[43][45], Harray[44][45], Harray[45][45], Harray[46][45], Harray[47][45], Harray[48][45], Harray[49][45], Harray[50][45], Harray[51][45], Harray[52][45], Harray[53][45], Harray[54][45], Harray[55][45], Harray[56][45], Harray[57][45], Harray[58][45], Harray[59][45], Harray[60][45], Harray[61][45], Harray[62][45], Harray[63][45], Harray[64][45], Harray[65][45], Harray[66][45], Harray[67][45], Harray[68][45], Harray[69][45], Harray[70][45], Harray[71][45], Harray[72][45], Harray[73][45], Harray[74][45], Harray[75][45], Harray[76][45], Harray[77][45], Harray[78][45], Harray[79][45], Harray[80][45], Harray[81][45], Harray[82][45], Harray[83][45], Harray[84][45], Harray[85][45], Harray[86][45], Harray[87][45], Harray[88][45], Harray[89][45], Harray[90][45], Harray[91][45], Harray[92][45], Harray[93][45], Harray[94][45], Harray[95][45], Harray[96][45], Harray[97][45], Harray[98][45], Harray[99][45], Harray[100][45], Harray[101][45], Harray[102][45], Harray[103][45], Harray[104][45], Harray[105][45], Harray[106][45], Harray[107][45], Harray[108][45], Harray[109][45], Harray[110][45], Harray[111][45], Harray[112][45], Harray[113][45], Harray[114][45], Harray[115][45], Harray[116][45], Harray[117][45], Harray[118][45], Harray[119][45], Harray[120][45], Harray[121][45], Harray[122][45], Harray[123][45], Harray[124][45], Harray[125][45], Harray[126][45], Harray[127][45]};
assign h_col_46 = {Harray[0][46], Harray[1][46], Harray[2][46], Harray[3][46], Harray[4][46], Harray[5][46], Harray[6][46], Harray[7][46], Harray[8][46], Harray[9][46], Harray[10][46], Harray[11][46], Harray[12][46], Harray[13][46], Harray[14][46], Harray[15][46], Harray[16][46], Harray[17][46], Harray[18][46], Harray[19][46], Harray[20][46], Harray[21][46], Harray[22][46], Harray[23][46], Harray[24][46], Harray[25][46], Harray[26][46], Harray[27][46], Harray[28][46], Harray[29][46], Harray[30][46], Harray[31][46], Harray[32][46], Harray[33][46], Harray[34][46], Harray[35][46], Harray[36][46], Harray[37][46], Harray[38][46], Harray[39][46], Harray[40][46], Harray[41][46], Harray[42][46], Harray[43][46], Harray[44][46], Harray[45][46], Harray[46][46], Harray[47][46], Harray[48][46], Harray[49][46], Harray[50][46], Harray[51][46], Harray[52][46], Harray[53][46], Harray[54][46], Harray[55][46], Harray[56][46], Harray[57][46], Harray[58][46], Harray[59][46], Harray[60][46], Harray[61][46], Harray[62][46], Harray[63][46], Harray[64][46], Harray[65][46], Harray[66][46], Harray[67][46], Harray[68][46], Harray[69][46], Harray[70][46], Harray[71][46], Harray[72][46], Harray[73][46], Harray[74][46], Harray[75][46], Harray[76][46], Harray[77][46], Harray[78][46], Harray[79][46], Harray[80][46], Harray[81][46], Harray[82][46], Harray[83][46], Harray[84][46], Harray[85][46], Harray[86][46], Harray[87][46], Harray[88][46], Harray[89][46], Harray[90][46], Harray[91][46], Harray[92][46], Harray[93][46], Harray[94][46], Harray[95][46], Harray[96][46], Harray[97][46], Harray[98][46], Harray[99][46], Harray[100][46], Harray[101][46], Harray[102][46], Harray[103][46], Harray[104][46], Harray[105][46], Harray[106][46], Harray[107][46], Harray[108][46], Harray[109][46], Harray[110][46], Harray[111][46], Harray[112][46], Harray[113][46], Harray[114][46], Harray[115][46], Harray[116][46], Harray[117][46], Harray[118][46], Harray[119][46], Harray[120][46], Harray[121][46], Harray[122][46], Harray[123][46], Harray[124][46], Harray[125][46], Harray[126][46], Harray[127][46]};
assign h_col_47 = {Harray[0][47], Harray[1][47], Harray[2][47], Harray[3][47], Harray[4][47], Harray[5][47], Harray[6][47], Harray[7][47], Harray[8][47], Harray[9][47], Harray[10][47], Harray[11][47], Harray[12][47], Harray[13][47], Harray[14][47], Harray[15][47], Harray[16][47], Harray[17][47], Harray[18][47], Harray[19][47], Harray[20][47], Harray[21][47], Harray[22][47], Harray[23][47], Harray[24][47], Harray[25][47], Harray[26][47], Harray[27][47], Harray[28][47], Harray[29][47], Harray[30][47], Harray[31][47], Harray[32][47], Harray[33][47], Harray[34][47], Harray[35][47], Harray[36][47], Harray[37][47], Harray[38][47], Harray[39][47], Harray[40][47], Harray[41][47], Harray[42][47], Harray[43][47], Harray[44][47], Harray[45][47], Harray[46][47], Harray[47][47], Harray[48][47], Harray[49][47], Harray[50][47], Harray[51][47], Harray[52][47], Harray[53][47], Harray[54][47], Harray[55][47], Harray[56][47], Harray[57][47], Harray[58][47], Harray[59][47], Harray[60][47], Harray[61][47], Harray[62][47], Harray[63][47], Harray[64][47], Harray[65][47], Harray[66][47], Harray[67][47], Harray[68][47], Harray[69][47], Harray[70][47], Harray[71][47], Harray[72][47], Harray[73][47], Harray[74][47], Harray[75][47], Harray[76][47], Harray[77][47], Harray[78][47], Harray[79][47], Harray[80][47], Harray[81][47], Harray[82][47], Harray[83][47], Harray[84][47], Harray[85][47], Harray[86][47], Harray[87][47], Harray[88][47], Harray[89][47], Harray[90][47], Harray[91][47], Harray[92][47], Harray[93][47], Harray[94][47], Harray[95][47], Harray[96][47], Harray[97][47], Harray[98][47], Harray[99][47], Harray[100][47], Harray[101][47], Harray[102][47], Harray[103][47], Harray[104][47], Harray[105][47], Harray[106][47], Harray[107][47], Harray[108][47], Harray[109][47], Harray[110][47], Harray[111][47], Harray[112][47], Harray[113][47], Harray[114][47], Harray[115][47], Harray[116][47], Harray[117][47], Harray[118][47], Harray[119][47], Harray[120][47], Harray[121][47], Harray[122][47], Harray[123][47], Harray[124][47], Harray[125][47], Harray[126][47], Harray[127][47]};
assign h_col_48 = {Harray[0][48], Harray[1][48], Harray[2][48], Harray[3][48], Harray[4][48], Harray[5][48], Harray[6][48], Harray[7][48], Harray[8][48], Harray[9][48], Harray[10][48], Harray[11][48], Harray[12][48], Harray[13][48], Harray[14][48], Harray[15][48], Harray[16][48], Harray[17][48], Harray[18][48], Harray[19][48], Harray[20][48], Harray[21][48], Harray[22][48], Harray[23][48], Harray[24][48], Harray[25][48], Harray[26][48], Harray[27][48], Harray[28][48], Harray[29][48], Harray[30][48], Harray[31][48], Harray[32][48], Harray[33][48], Harray[34][48], Harray[35][48], Harray[36][48], Harray[37][48], Harray[38][48], Harray[39][48], Harray[40][48], Harray[41][48], Harray[42][48], Harray[43][48], Harray[44][48], Harray[45][48], Harray[46][48], Harray[47][48], Harray[48][48], Harray[49][48], Harray[50][48], Harray[51][48], Harray[52][48], Harray[53][48], Harray[54][48], Harray[55][48], Harray[56][48], Harray[57][48], Harray[58][48], Harray[59][48], Harray[60][48], Harray[61][48], Harray[62][48], Harray[63][48], Harray[64][48], Harray[65][48], Harray[66][48], Harray[67][48], Harray[68][48], Harray[69][48], Harray[70][48], Harray[71][48], Harray[72][48], Harray[73][48], Harray[74][48], Harray[75][48], Harray[76][48], Harray[77][48], Harray[78][48], Harray[79][48], Harray[80][48], Harray[81][48], Harray[82][48], Harray[83][48], Harray[84][48], Harray[85][48], Harray[86][48], Harray[87][48], Harray[88][48], Harray[89][48], Harray[90][48], Harray[91][48], Harray[92][48], Harray[93][48], Harray[94][48], Harray[95][48], Harray[96][48], Harray[97][48], Harray[98][48], Harray[99][48], Harray[100][48], Harray[101][48], Harray[102][48], Harray[103][48], Harray[104][48], Harray[105][48], Harray[106][48], Harray[107][48], Harray[108][48], Harray[109][48], Harray[110][48], Harray[111][48], Harray[112][48], Harray[113][48], Harray[114][48], Harray[115][48], Harray[116][48], Harray[117][48], Harray[118][48], Harray[119][48], Harray[120][48], Harray[121][48], Harray[122][48], Harray[123][48], Harray[124][48], Harray[125][48], Harray[126][48], Harray[127][48]};
assign h_col_49 = {Harray[0][49], Harray[1][49], Harray[2][49], Harray[3][49], Harray[4][49], Harray[5][49], Harray[6][49], Harray[7][49], Harray[8][49], Harray[9][49], Harray[10][49], Harray[11][49], Harray[12][49], Harray[13][49], Harray[14][49], Harray[15][49], Harray[16][49], Harray[17][49], Harray[18][49], Harray[19][49], Harray[20][49], Harray[21][49], Harray[22][49], Harray[23][49], Harray[24][49], Harray[25][49], Harray[26][49], Harray[27][49], Harray[28][49], Harray[29][49], Harray[30][49], Harray[31][49], Harray[32][49], Harray[33][49], Harray[34][49], Harray[35][49], Harray[36][49], Harray[37][49], Harray[38][49], Harray[39][49], Harray[40][49], Harray[41][49], Harray[42][49], Harray[43][49], Harray[44][49], Harray[45][49], Harray[46][49], Harray[47][49], Harray[48][49], Harray[49][49], Harray[50][49], Harray[51][49], Harray[52][49], Harray[53][49], Harray[54][49], Harray[55][49], Harray[56][49], Harray[57][49], Harray[58][49], Harray[59][49], Harray[60][49], Harray[61][49], Harray[62][49], Harray[63][49], Harray[64][49], Harray[65][49], Harray[66][49], Harray[67][49], Harray[68][49], Harray[69][49], Harray[70][49], Harray[71][49], Harray[72][49], Harray[73][49], Harray[74][49], Harray[75][49], Harray[76][49], Harray[77][49], Harray[78][49], Harray[79][49], Harray[80][49], Harray[81][49], Harray[82][49], Harray[83][49], Harray[84][49], Harray[85][49], Harray[86][49], Harray[87][49], Harray[88][49], Harray[89][49], Harray[90][49], Harray[91][49], Harray[92][49], Harray[93][49], Harray[94][49], Harray[95][49], Harray[96][49], Harray[97][49], Harray[98][49], Harray[99][49], Harray[100][49], Harray[101][49], Harray[102][49], Harray[103][49], Harray[104][49], Harray[105][49], Harray[106][49], Harray[107][49], Harray[108][49], Harray[109][49], Harray[110][49], Harray[111][49], Harray[112][49], Harray[113][49], Harray[114][49], Harray[115][49], Harray[116][49], Harray[117][49], Harray[118][49], Harray[119][49], Harray[120][49], Harray[121][49], Harray[122][49], Harray[123][49], Harray[124][49], Harray[125][49], Harray[126][49], Harray[127][49]};
assign h_col_50 = {Harray[0][50], Harray[1][50], Harray[2][50], Harray[3][50], Harray[4][50], Harray[5][50], Harray[6][50], Harray[7][50], Harray[8][50], Harray[9][50], Harray[10][50], Harray[11][50], Harray[12][50], Harray[13][50], Harray[14][50], Harray[15][50], Harray[16][50], Harray[17][50], Harray[18][50], Harray[19][50], Harray[20][50], Harray[21][50], Harray[22][50], Harray[23][50], Harray[24][50], Harray[25][50], Harray[26][50], Harray[27][50], Harray[28][50], Harray[29][50], Harray[30][50], Harray[31][50], Harray[32][50], Harray[33][50], Harray[34][50], Harray[35][50], Harray[36][50], Harray[37][50], Harray[38][50], Harray[39][50], Harray[40][50], Harray[41][50], Harray[42][50], Harray[43][50], Harray[44][50], Harray[45][50], Harray[46][50], Harray[47][50], Harray[48][50], Harray[49][50], Harray[50][50], Harray[51][50], Harray[52][50], Harray[53][50], Harray[54][50], Harray[55][50], Harray[56][50], Harray[57][50], Harray[58][50], Harray[59][50], Harray[60][50], Harray[61][50], Harray[62][50], Harray[63][50], Harray[64][50], Harray[65][50], Harray[66][50], Harray[67][50], Harray[68][50], Harray[69][50], Harray[70][50], Harray[71][50], Harray[72][50], Harray[73][50], Harray[74][50], Harray[75][50], Harray[76][50], Harray[77][50], Harray[78][50], Harray[79][50], Harray[80][50], Harray[81][50], Harray[82][50], Harray[83][50], Harray[84][50], Harray[85][50], Harray[86][50], Harray[87][50], Harray[88][50], Harray[89][50], Harray[90][50], Harray[91][50], Harray[92][50], Harray[93][50], Harray[94][50], Harray[95][50], Harray[96][50], Harray[97][50], Harray[98][50], Harray[99][50], Harray[100][50], Harray[101][50], Harray[102][50], Harray[103][50], Harray[104][50], Harray[105][50], Harray[106][50], Harray[107][50], Harray[108][50], Harray[109][50], Harray[110][50], Harray[111][50], Harray[112][50], Harray[113][50], Harray[114][50], Harray[115][50], Harray[116][50], Harray[117][50], Harray[118][50], Harray[119][50], Harray[120][50], Harray[121][50], Harray[122][50], Harray[123][50], Harray[124][50], Harray[125][50], Harray[126][50], Harray[127][50]};
assign h_col_51 = {Harray[0][51], Harray[1][51], Harray[2][51], Harray[3][51], Harray[4][51], Harray[5][51], Harray[6][51], Harray[7][51], Harray[8][51], Harray[9][51], Harray[10][51], Harray[11][51], Harray[12][51], Harray[13][51], Harray[14][51], Harray[15][51], Harray[16][51], Harray[17][51], Harray[18][51], Harray[19][51], Harray[20][51], Harray[21][51], Harray[22][51], Harray[23][51], Harray[24][51], Harray[25][51], Harray[26][51], Harray[27][51], Harray[28][51], Harray[29][51], Harray[30][51], Harray[31][51], Harray[32][51], Harray[33][51], Harray[34][51], Harray[35][51], Harray[36][51], Harray[37][51], Harray[38][51], Harray[39][51], Harray[40][51], Harray[41][51], Harray[42][51], Harray[43][51], Harray[44][51], Harray[45][51], Harray[46][51], Harray[47][51], Harray[48][51], Harray[49][51], Harray[50][51], Harray[51][51], Harray[52][51], Harray[53][51], Harray[54][51], Harray[55][51], Harray[56][51], Harray[57][51], Harray[58][51], Harray[59][51], Harray[60][51], Harray[61][51], Harray[62][51], Harray[63][51], Harray[64][51], Harray[65][51], Harray[66][51], Harray[67][51], Harray[68][51], Harray[69][51], Harray[70][51], Harray[71][51], Harray[72][51], Harray[73][51], Harray[74][51], Harray[75][51], Harray[76][51], Harray[77][51], Harray[78][51], Harray[79][51], Harray[80][51], Harray[81][51], Harray[82][51], Harray[83][51], Harray[84][51], Harray[85][51], Harray[86][51], Harray[87][51], Harray[88][51], Harray[89][51], Harray[90][51], Harray[91][51], Harray[92][51], Harray[93][51], Harray[94][51], Harray[95][51], Harray[96][51], Harray[97][51], Harray[98][51], Harray[99][51], Harray[100][51], Harray[101][51], Harray[102][51], Harray[103][51], Harray[104][51], Harray[105][51], Harray[106][51], Harray[107][51], Harray[108][51], Harray[109][51], Harray[110][51], Harray[111][51], Harray[112][51], Harray[113][51], Harray[114][51], Harray[115][51], Harray[116][51], Harray[117][51], Harray[118][51], Harray[119][51], Harray[120][51], Harray[121][51], Harray[122][51], Harray[123][51], Harray[124][51], Harray[125][51], Harray[126][51], Harray[127][51]};
assign h_col_52 = {Harray[0][52], Harray[1][52], Harray[2][52], Harray[3][52], Harray[4][52], Harray[5][52], Harray[6][52], Harray[7][52], Harray[8][52], Harray[9][52], Harray[10][52], Harray[11][52], Harray[12][52], Harray[13][52], Harray[14][52], Harray[15][52], Harray[16][52], Harray[17][52], Harray[18][52], Harray[19][52], Harray[20][52], Harray[21][52], Harray[22][52], Harray[23][52], Harray[24][52], Harray[25][52], Harray[26][52], Harray[27][52], Harray[28][52], Harray[29][52], Harray[30][52], Harray[31][52], Harray[32][52], Harray[33][52], Harray[34][52], Harray[35][52], Harray[36][52], Harray[37][52], Harray[38][52], Harray[39][52], Harray[40][52], Harray[41][52], Harray[42][52], Harray[43][52], Harray[44][52], Harray[45][52], Harray[46][52], Harray[47][52], Harray[48][52], Harray[49][52], Harray[50][52], Harray[51][52], Harray[52][52], Harray[53][52], Harray[54][52], Harray[55][52], Harray[56][52], Harray[57][52], Harray[58][52], Harray[59][52], Harray[60][52], Harray[61][52], Harray[62][52], Harray[63][52], Harray[64][52], Harray[65][52], Harray[66][52], Harray[67][52], Harray[68][52], Harray[69][52], Harray[70][52], Harray[71][52], Harray[72][52], Harray[73][52], Harray[74][52], Harray[75][52], Harray[76][52], Harray[77][52], Harray[78][52], Harray[79][52], Harray[80][52], Harray[81][52], Harray[82][52], Harray[83][52], Harray[84][52], Harray[85][52], Harray[86][52], Harray[87][52], Harray[88][52], Harray[89][52], Harray[90][52], Harray[91][52], Harray[92][52], Harray[93][52], Harray[94][52], Harray[95][52], Harray[96][52], Harray[97][52], Harray[98][52], Harray[99][52], Harray[100][52], Harray[101][52], Harray[102][52], Harray[103][52], Harray[104][52], Harray[105][52], Harray[106][52], Harray[107][52], Harray[108][52], Harray[109][52], Harray[110][52], Harray[111][52], Harray[112][52], Harray[113][52], Harray[114][52], Harray[115][52], Harray[116][52], Harray[117][52], Harray[118][52], Harray[119][52], Harray[120][52], Harray[121][52], Harray[122][52], Harray[123][52], Harray[124][52], Harray[125][52], Harray[126][52], Harray[127][52]};
assign h_col_53 = {Harray[0][53], Harray[1][53], Harray[2][53], Harray[3][53], Harray[4][53], Harray[5][53], Harray[6][53], Harray[7][53], Harray[8][53], Harray[9][53], Harray[10][53], Harray[11][53], Harray[12][53], Harray[13][53], Harray[14][53], Harray[15][53], Harray[16][53], Harray[17][53], Harray[18][53], Harray[19][53], Harray[20][53], Harray[21][53], Harray[22][53], Harray[23][53], Harray[24][53], Harray[25][53], Harray[26][53], Harray[27][53], Harray[28][53], Harray[29][53], Harray[30][53], Harray[31][53], Harray[32][53], Harray[33][53], Harray[34][53], Harray[35][53], Harray[36][53], Harray[37][53], Harray[38][53], Harray[39][53], Harray[40][53], Harray[41][53], Harray[42][53], Harray[43][53], Harray[44][53], Harray[45][53], Harray[46][53], Harray[47][53], Harray[48][53], Harray[49][53], Harray[50][53], Harray[51][53], Harray[52][53], Harray[53][53], Harray[54][53], Harray[55][53], Harray[56][53], Harray[57][53], Harray[58][53], Harray[59][53], Harray[60][53], Harray[61][53], Harray[62][53], Harray[63][53], Harray[64][53], Harray[65][53], Harray[66][53], Harray[67][53], Harray[68][53], Harray[69][53], Harray[70][53], Harray[71][53], Harray[72][53], Harray[73][53], Harray[74][53], Harray[75][53], Harray[76][53], Harray[77][53], Harray[78][53], Harray[79][53], Harray[80][53], Harray[81][53], Harray[82][53], Harray[83][53], Harray[84][53], Harray[85][53], Harray[86][53], Harray[87][53], Harray[88][53], Harray[89][53], Harray[90][53], Harray[91][53], Harray[92][53], Harray[93][53], Harray[94][53], Harray[95][53], Harray[96][53], Harray[97][53], Harray[98][53], Harray[99][53], Harray[100][53], Harray[101][53], Harray[102][53], Harray[103][53], Harray[104][53], Harray[105][53], Harray[106][53], Harray[107][53], Harray[108][53], Harray[109][53], Harray[110][53], Harray[111][53], Harray[112][53], Harray[113][53], Harray[114][53], Harray[115][53], Harray[116][53], Harray[117][53], Harray[118][53], Harray[119][53], Harray[120][53], Harray[121][53], Harray[122][53], Harray[123][53], Harray[124][53], Harray[125][53], Harray[126][53], Harray[127][53]};
assign h_col_54 = {Harray[0][54], Harray[1][54], Harray[2][54], Harray[3][54], Harray[4][54], Harray[5][54], Harray[6][54], Harray[7][54], Harray[8][54], Harray[9][54], Harray[10][54], Harray[11][54], Harray[12][54], Harray[13][54], Harray[14][54], Harray[15][54], Harray[16][54], Harray[17][54], Harray[18][54], Harray[19][54], Harray[20][54], Harray[21][54], Harray[22][54], Harray[23][54], Harray[24][54], Harray[25][54], Harray[26][54], Harray[27][54], Harray[28][54], Harray[29][54], Harray[30][54], Harray[31][54], Harray[32][54], Harray[33][54], Harray[34][54], Harray[35][54], Harray[36][54], Harray[37][54], Harray[38][54], Harray[39][54], Harray[40][54], Harray[41][54], Harray[42][54], Harray[43][54], Harray[44][54], Harray[45][54], Harray[46][54], Harray[47][54], Harray[48][54], Harray[49][54], Harray[50][54], Harray[51][54], Harray[52][54], Harray[53][54], Harray[54][54], Harray[55][54], Harray[56][54], Harray[57][54], Harray[58][54], Harray[59][54], Harray[60][54], Harray[61][54], Harray[62][54], Harray[63][54], Harray[64][54], Harray[65][54], Harray[66][54], Harray[67][54], Harray[68][54], Harray[69][54], Harray[70][54], Harray[71][54], Harray[72][54], Harray[73][54], Harray[74][54], Harray[75][54], Harray[76][54], Harray[77][54], Harray[78][54], Harray[79][54], Harray[80][54], Harray[81][54], Harray[82][54], Harray[83][54], Harray[84][54], Harray[85][54], Harray[86][54], Harray[87][54], Harray[88][54], Harray[89][54], Harray[90][54], Harray[91][54], Harray[92][54], Harray[93][54], Harray[94][54], Harray[95][54], Harray[96][54], Harray[97][54], Harray[98][54], Harray[99][54], Harray[100][54], Harray[101][54], Harray[102][54], Harray[103][54], Harray[104][54], Harray[105][54], Harray[106][54], Harray[107][54], Harray[108][54], Harray[109][54], Harray[110][54], Harray[111][54], Harray[112][54], Harray[113][54], Harray[114][54], Harray[115][54], Harray[116][54], Harray[117][54], Harray[118][54], Harray[119][54], Harray[120][54], Harray[121][54], Harray[122][54], Harray[123][54], Harray[124][54], Harray[125][54], Harray[126][54], Harray[127][54]};
assign h_col_55 = {Harray[0][55], Harray[1][55], Harray[2][55], Harray[3][55], Harray[4][55], Harray[5][55], Harray[6][55], Harray[7][55], Harray[8][55], Harray[9][55], Harray[10][55], Harray[11][55], Harray[12][55], Harray[13][55], Harray[14][55], Harray[15][55], Harray[16][55], Harray[17][55], Harray[18][55], Harray[19][55], Harray[20][55], Harray[21][55], Harray[22][55], Harray[23][55], Harray[24][55], Harray[25][55], Harray[26][55], Harray[27][55], Harray[28][55], Harray[29][55], Harray[30][55], Harray[31][55], Harray[32][55], Harray[33][55], Harray[34][55], Harray[35][55], Harray[36][55], Harray[37][55], Harray[38][55], Harray[39][55], Harray[40][55], Harray[41][55], Harray[42][55], Harray[43][55], Harray[44][55], Harray[45][55], Harray[46][55], Harray[47][55], Harray[48][55], Harray[49][55], Harray[50][55], Harray[51][55], Harray[52][55], Harray[53][55], Harray[54][55], Harray[55][55], Harray[56][55], Harray[57][55], Harray[58][55], Harray[59][55], Harray[60][55], Harray[61][55], Harray[62][55], Harray[63][55], Harray[64][55], Harray[65][55], Harray[66][55], Harray[67][55], Harray[68][55], Harray[69][55], Harray[70][55], Harray[71][55], Harray[72][55], Harray[73][55], Harray[74][55], Harray[75][55], Harray[76][55], Harray[77][55], Harray[78][55], Harray[79][55], Harray[80][55], Harray[81][55], Harray[82][55], Harray[83][55], Harray[84][55], Harray[85][55], Harray[86][55], Harray[87][55], Harray[88][55], Harray[89][55], Harray[90][55], Harray[91][55], Harray[92][55], Harray[93][55], Harray[94][55], Harray[95][55], Harray[96][55], Harray[97][55], Harray[98][55], Harray[99][55], Harray[100][55], Harray[101][55], Harray[102][55], Harray[103][55], Harray[104][55], Harray[105][55], Harray[106][55], Harray[107][55], Harray[108][55], Harray[109][55], Harray[110][55], Harray[111][55], Harray[112][55], Harray[113][55], Harray[114][55], Harray[115][55], Harray[116][55], Harray[117][55], Harray[118][55], Harray[119][55], Harray[120][55], Harray[121][55], Harray[122][55], Harray[123][55], Harray[124][55], Harray[125][55], Harray[126][55], Harray[127][55]};
assign h_col_56 = {Harray[0][56], Harray[1][56], Harray[2][56], Harray[3][56], Harray[4][56], Harray[5][56], Harray[6][56], Harray[7][56], Harray[8][56], Harray[9][56], Harray[10][56], Harray[11][56], Harray[12][56], Harray[13][56], Harray[14][56], Harray[15][56], Harray[16][56], Harray[17][56], Harray[18][56], Harray[19][56], Harray[20][56], Harray[21][56], Harray[22][56], Harray[23][56], Harray[24][56], Harray[25][56], Harray[26][56], Harray[27][56], Harray[28][56], Harray[29][56], Harray[30][56], Harray[31][56], Harray[32][56], Harray[33][56], Harray[34][56], Harray[35][56], Harray[36][56], Harray[37][56], Harray[38][56], Harray[39][56], Harray[40][56], Harray[41][56], Harray[42][56], Harray[43][56], Harray[44][56], Harray[45][56], Harray[46][56], Harray[47][56], Harray[48][56], Harray[49][56], Harray[50][56], Harray[51][56], Harray[52][56], Harray[53][56], Harray[54][56], Harray[55][56], Harray[56][56], Harray[57][56], Harray[58][56], Harray[59][56], Harray[60][56], Harray[61][56], Harray[62][56], Harray[63][56], Harray[64][56], Harray[65][56], Harray[66][56], Harray[67][56], Harray[68][56], Harray[69][56], Harray[70][56], Harray[71][56], Harray[72][56], Harray[73][56], Harray[74][56], Harray[75][56], Harray[76][56], Harray[77][56], Harray[78][56], Harray[79][56], Harray[80][56], Harray[81][56], Harray[82][56], Harray[83][56], Harray[84][56], Harray[85][56], Harray[86][56], Harray[87][56], Harray[88][56], Harray[89][56], Harray[90][56], Harray[91][56], Harray[92][56], Harray[93][56], Harray[94][56], Harray[95][56], Harray[96][56], Harray[97][56], Harray[98][56], Harray[99][56], Harray[100][56], Harray[101][56], Harray[102][56], Harray[103][56], Harray[104][56], Harray[105][56], Harray[106][56], Harray[107][56], Harray[108][56], Harray[109][56], Harray[110][56], Harray[111][56], Harray[112][56], Harray[113][56], Harray[114][56], Harray[115][56], Harray[116][56], Harray[117][56], Harray[118][56], Harray[119][56], Harray[120][56], Harray[121][56], Harray[122][56], Harray[123][56], Harray[124][56], Harray[125][56], Harray[126][56], Harray[127][56]};
assign h_col_57 = {Harray[0][57], Harray[1][57], Harray[2][57], Harray[3][57], Harray[4][57], Harray[5][57], Harray[6][57], Harray[7][57], Harray[8][57], Harray[9][57], Harray[10][57], Harray[11][57], Harray[12][57], Harray[13][57], Harray[14][57], Harray[15][57], Harray[16][57], Harray[17][57], Harray[18][57], Harray[19][57], Harray[20][57], Harray[21][57], Harray[22][57], Harray[23][57], Harray[24][57], Harray[25][57], Harray[26][57], Harray[27][57], Harray[28][57], Harray[29][57], Harray[30][57], Harray[31][57], Harray[32][57], Harray[33][57], Harray[34][57], Harray[35][57], Harray[36][57], Harray[37][57], Harray[38][57], Harray[39][57], Harray[40][57], Harray[41][57], Harray[42][57], Harray[43][57], Harray[44][57], Harray[45][57], Harray[46][57], Harray[47][57], Harray[48][57], Harray[49][57], Harray[50][57], Harray[51][57], Harray[52][57], Harray[53][57], Harray[54][57], Harray[55][57], Harray[56][57], Harray[57][57], Harray[58][57], Harray[59][57], Harray[60][57], Harray[61][57], Harray[62][57], Harray[63][57], Harray[64][57], Harray[65][57], Harray[66][57], Harray[67][57], Harray[68][57], Harray[69][57], Harray[70][57], Harray[71][57], Harray[72][57], Harray[73][57], Harray[74][57], Harray[75][57], Harray[76][57], Harray[77][57], Harray[78][57], Harray[79][57], Harray[80][57], Harray[81][57], Harray[82][57], Harray[83][57], Harray[84][57], Harray[85][57], Harray[86][57], Harray[87][57], Harray[88][57], Harray[89][57], Harray[90][57], Harray[91][57], Harray[92][57], Harray[93][57], Harray[94][57], Harray[95][57], Harray[96][57], Harray[97][57], Harray[98][57], Harray[99][57], Harray[100][57], Harray[101][57], Harray[102][57], Harray[103][57], Harray[104][57], Harray[105][57], Harray[106][57], Harray[107][57], Harray[108][57], Harray[109][57], Harray[110][57], Harray[111][57], Harray[112][57], Harray[113][57], Harray[114][57], Harray[115][57], Harray[116][57], Harray[117][57], Harray[118][57], Harray[119][57], Harray[120][57], Harray[121][57], Harray[122][57], Harray[123][57], Harray[124][57], Harray[125][57], Harray[126][57], Harray[127][57]};
assign h_col_58 = {Harray[0][58], Harray[1][58], Harray[2][58], Harray[3][58], Harray[4][58], Harray[5][58], Harray[6][58], Harray[7][58], Harray[8][58], Harray[9][58], Harray[10][58], Harray[11][58], Harray[12][58], Harray[13][58], Harray[14][58], Harray[15][58], Harray[16][58], Harray[17][58], Harray[18][58], Harray[19][58], Harray[20][58], Harray[21][58], Harray[22][58], Harray[23][58], Harray[24][58], Harray[25][58], Harray[26][58], Harray[27][58], Harray[28][58], Harray[29][58], Harray[30][58], Harray[31][58], Harray[32][58], Harray[33][58], Harray[34][58], Harray[35][58], Harray[36][58], Harray[37][58], Harray[38][58], Harray[39][58], Harray[40][58], Harray[41][58], Harray[42][58], Harray[43][58], Harray[44][58], Harray[45][58], Harray[46][58], Harray[47][58], Harray[48][58], Harray[49][58], Harray[50][58], Harray[51][58], Harray[52][58], Harray[53][58], Harray[54][58], Harray[55][58], Harray[56][58], Harray[57][58], Harray[58][58], Harray[59][58], Harray[60][58], Harray[61][58], Harray[62][58], Harray[63][58], Harray[64][58], Harray[65][58], Harray[66][58], Harray[67][58], Harray[68][58], Harray[69][58], Harray[70][58], Harray[71][58], Harray[72][58], Harray[73][58], Harray[74][58], Harray[75][58], Harray[76][58], Harray[77][58], Harray[78][58], Harray[79][58], Harray[80][58], Harray[81][58], Harray[82][58], Harray[83][58], Harray[84][58], Harray[85][58], Harray[86][58], Harray[87][58], Harray[88][58], Harray[89][58], Harray[90][58], Harray[91][58], Harray[92][58], Harray[93][58], Harray[94][58], Harray[95][58], Harray[96][58], Harray[97][58], Harray[98][58], Harray[99][58], Harray[100][58], Harray[101][58], Harray[102][58], Harray[103][58], Harray[104][58], Harray[105][58], Harray[106][58], Harray[107][58], Harray[108][58], Harray[109][58], Harray[110][58], Harray[111][58], Harray[112][58], Harray[113][58], Harray[114][58], Harray[115][58], Harray[116][58], Harray[117][58], Harray[118][58], Harray[119][58], Harray[120][58], Harray[121][58], Harray[122][58], Harray[123][58], Harray[124][58], Harray[125][58], Harray[126][58], Harray[127][58]};
assign h_col_59 = {Harray[0][59], Harray[1][59], Harray[2][59], Harray[3][59], Harray[4][59], Harray[5][59], Harray[6][59], Harray[7][59], Harray[8][59], Harray[9][59], Harray[10][59], Harray[11][59], Harray[12][59], Harray[13][59], Harray[14][59], Harray[15][59], Harray[16][59], Harray[17][59], Harray[18][59], Harray[19][59], Harray[20][59], Harray[21][59], Harray[22][59], Harray[23][59], Harray[24][59], Harray[25][59], Harray[26][59], Harray[27][59], Harray[28][59], Harray[29][59], Harray[30][59], Harray[31][59], Harray[32][59], Harray[33][59], Harray[34][59], Harray[35][59], Harray[36][59], Harray[37][59], Harray[38][59], Harray[39][59], Harray[40][59], Harray[41][59], Harray[42][59], Harray[43][59], Harray[44][59], Harray[45][59], Harray[46][59], Harray[47][59], Harray[48][59], Harray[49][59], Harray[50][59], Harray[51][59], Harray[52][59], Harray[53][59], Harray[54][59], Harray[55][59], Harray[56][59], Harray[57][59], Harray[58][59], Harray[59][59], Harray[60][59], Harray[61][59], Harray[62][59], Harray[63][59], Harray[64][59], Harray[65][59], Harray[66][59], Harray[67][59], Harray[68][59], Harray[69][59], Harray[70][59], Harray[71][59], Harray[72][59], Harray[73][59], Harray[74][59], Harray[75][59], Harray[76][59], Harray[77][59], Harray[78][59], Harray[79][59], Harray[80][59], Harray[81][59], Harray[82][59], Harray[83][59], Harray[84][59], Harray[85][59], Harray[86][59], Harray[87][59], Harray[88][59], Harray[89][59], Harray[90][59], Harray[91][59], Harray[92][59], Harray[93][59], Harray[94][59], Harray[95][59], Harray[96][59], Harray[97][59], Harray[98][59], Harray[99][59], Harray[100][59], Harray[101][59], Harray[102][59], Harray[103][59], Harray[104][59], Harray[105][59], Harray[106][59], Harray[107][59], Harray[108][59], Harray[109][59], Harray[110][59], Harray[111][59], Harray[112][59], Harray[113][59], Harray[114][59], Harray[115][59], Harray[116][59], Harray[117][59], Harray[118][59], Harray[119][59], Harray[120][59], Harray[121][59], Harray[122][59], Harray[123][59], Harray[124][59], Harray[125][59], Harray[126][59], Harray[127][59]};
assign h_col_60 = {Harray[0][60], Harray[1][60], Harray[2][60], Harray[3][60], Harray[4][60], Harray[5][60], Harray[6][60], Harray[7][60], Harray[8][60], Harray[9][60], Harray[10][60], Harray[11][60], Harray[12][60], Harray[13][60], Harray[14][60], Harray[15][60], Harray[16][60], Harray[17][60], Harray[18][60], Harray[19][60], Harray[20][60], Harray[21][60], Harray[22][60], Harray[23][60], Harray[24][60], Harray[25][60], Harray[26][60], Harray[27][60], Harray[28][60], Harray[29][60], Harray[30][60], Harray[31][60], Harray[32][60], Harray[33][60], Harray[34][60], Harray[35][60], Harray[36][60], Harray[37][60], Harray[38][60], Harray[39][60], Harray[40][60], Harray[41][60], Harray[42][60], Harray[43][60], Harray[44][60], Harray[45][60], Harray[46][60], Harray[47][60], Harray[48][60], Harray[49][60], Harray[50][60], Harray[51][60], Harray[52][60], Harray[53][60], Harray[54][60], Harray[55][60], Harray[56][60], Harray[57][60], Harray[58][60], Harray[59][60], Harray[60][60], Harray[61][60], Harray[62][60], Harray[63][60], Harray[64][60], Harray[65][60], Harray[66][60], Harray[67][60], Harray[68][60], Harray[69][60], Harray[70][60], Harray[71][60], Harray[72][60], Harray[73][60], Harray[74][60], Harray[75][60], Harray[76][60], Harray[77][60], Harray[78][60], Harray[79][60], Harray[80][60], Harray[81][60], Harray[82][60], Harray[83][60], Harray[84][60], Harray[85][60], Harray[86][60], Harray[87][60], Harray[88][60], Harray[89][60], Harray[90][60], Harray[91][60], Harray[92][60], Harray[93][60], Harray[94][60], Harray[95][60], Harray[96][60], Harray[97][60], Harray[98][60], Harray[99][60], Harray[100][60], Harray[101][60], Harray[102][60], Harray[103][60], Harray[104][60], Harray[105][60], Harray[106][60], Harray[107][60], Harray[108][60], Harray[109][60], Harray[110][60], Harray[111][60], Harray[112][60], Harray[113][60], Harray[114][60], Harray[115][60], Harray[116][60], Harray[117][60], Harray[118][60], Harray[119][60], Harray[120][60], Harray[121][60], Harray[122][60], Harray[123][60], Harray[124][60], Harray[125][60], Harray[126][60], Harray[127][60]};
assign h_col_61 = {Harray[0][61], Harray[1][61], Harray[2][61], Harray[3][61], Harray[4][61], Harray[5][61], Harray[6][61], Harray[7][61], Harray[8][61], Harray[9][61], Harray[10][61], Harray[11][61], Harray[12][61], Harray[13][61], Harray[14][61], Harray[15][61], Harray[16][61], Harray[17][61], Harray[18][61], Harray[19][61], Harray[20][61], Harray[21][61], Harray[22][61], Harray[23][61], Harray[24][61], Harray[25][61], Harray[26][61], Harray[27][61], Harray[28][61], Harray[29][61], Harray[30][61], Harray[31][61], Harray[32][61], Harray[33][61], Harray[34][61], Harray[35][61], Harray[36][61], Harray[37][61], Harray[38][61], Harray[39][61], Harray[40][61], Harray[41][61], Harray[42][61], Harray[43][61], Harray[44][61], Harray[45][61], Harray[46][61], Harray[47][61], Harray[48][61], Harray[49][61], Harray[50][61], Harray[51][61], Harray[52][61], Harray[53][61], Harray[54][61], Harray[55][61], Harray[56][61], Harray[57][61], Harray[58][61], Harray[59][61], Harray[60][61], Harray[61][61], Harray[62][61], Harray[63][61], Harray[64][61], Harray[65][61], Harray[66][61], Harray[67][61], Harray[68][61], Harray[69][61], Harray[70][61], Harray[71][61], Harray[72][61], Harray[73][61], Harray[74][61], Harray[75][61], Harray[76][61], Harray[77][61], Harray[78][61], Harray[79][61], Harray[80][61], Harray[81][61], Harray[82][61], Harray[83][61], Harray[84][61], Harray[85][61], Harray[86][61], Harray[87][61], Harray[88][61], Harray[89][61], Harray[90][61], Harray[91][61], Harray[92][61], Harray[93][61], Harray[94][61], Harray[95][61], Harray[96][61], Harray[97][61], Harray[98][61], Harray[99][61], Harray[100][61], Harray[101][61], Harray[102][61], Harray[103][61], Harray[104][61], Harray[105][61], Harray[106][61], Harray[107][61], Harray[108][61], Harray[109][61], Harray[110][61], Harray[111][61], Harray[112][61], Harray[113][61], Harray[114][61], Harray[115][61], Harray[116][61], Harray[117][61], Harray[118][61], Harray[119][61], Harray[120][61], Harray[121][61], Harray[122][61], Harray[123][61], Harray[124][61], Harray[125][61], Harray[126][61], Harray[127][61]};
assign h_col_62 = {Harray[0][62], Harray[1][62], Harray[2][62], Harray[3][62], Harray[4][62], Harray[5][62], Harray[6][62], Harray[7][62], Harray[8][62], Harray[9][62], Harray[10][62], Harray[11][62], Harray[12][62], Harray[13][62], Harray[14][62], Harray[15][62], Harray[16][62], Harray[17][62], Harray[18][62], Harray[19][62], Harray[20][62], Harray[21][62], Harray[22][62], Harray[23][62], Harray[24][62], Harray[25][62], Harray[26][62], Harray[27][62], Harray[28][62], Harray[29][62], Harray[30][62], Harray[31][62], Harray[32][62], Harray[33][62], Harray[34][62], Harray[35][62], Harray[36][62], Harray[37][62], Harray[38][62], Harray[39][62], Harray[40][62], Harray[41][62], Harray[42][62], Harray[43][62], Harray[44][62], Harray[45][62], Harray[46][62], Harray[47][62], Harray[48][62], Harray[49][62], Harray[50][62], Harray[51][62], Harray[52][62], Harray[53][62], Harray[54][62], Harray[55][62], Harray[56][62], Harray[57][62], Harray[58][62], Harray[59][62], Harray[60][62], Harray[61][62], Harray[62][62], Harray[63][62], Harray[64][62], Harray[65][62], Harray[66][62], Harray[67][62], Harray[68][62], Harray[69][62], Harray[70][62], Harray[71][62], Harray[72][62], Harray[73][62], Harray[74][62], Harray[75][62], Harray[76][62], Harray[77][62], Harray[78][62], Harray[79][62], Harray[80][62], Harray[81][62], Harray[82][62], Harray[83][62], Harray[84][62], Harray[85][62], Harray[86][62], Harray[87][62], Harray[88][62], Harray[89][62], Harray[90][62], Harray[91][62], Harray[92][62], Harray[93][62], Harray[94][62], Harray[95][62], Harray[96][62], Harray[97][62], Harray[98][62], Harray[99][62], Harray[100][62], Harray[101][62], Harray[102][62], Harray[103][62], Harray[104][62], Harray[105][62], Harray[106][62], Harray[107][62], Harray[108][62], Harray[109][62], Harray[110][62], Harray[111][62], Harray[112][62], Harray[113][62], Harray[114][62], Harray[115][62], Harray[116][62], Harray[117][62], Harray[118][62], Harray[119][62], Harray[120][62], Harray[121][62], Harray[122][62], Harray[123][62], Harray[124][62], Harray[125][62], Harray[126][62], Harray[127][62]};
assign h_col_63 = {Harray[0][63], Harray[1][63], Harray[2][63], Harray[3][63], Harray[4][63], Harray[5][63], Harray[6][63], Harray[7][63], Harray[8][63], Harray[9][63], Harray[10][63], Harray[11][63], Harray[12][63], Harray[13][63], Harray[14][63], Harray[15][63], Harray[16][63], Harray[17][63], Harray[18][63], Harray[19][63], Harray[20][63], Harray[21][63], Harray[22][63], Harray[23][63], Harray[24][63], Harray[25][63], Harray[26][63], Harray[27][63], Harray[28][63], Harray[29][63], Harray[30][63], Harray[31][63], Harray[32][63], Harray[33][63], Harray[34][63], Harray[35][63], Harray[36][63], Harray[37][63], Harray[38][63], Harray[39][63], Harray[40][63], Harray[41][63], Harray[42][63], Harray[43][63], Harray[44][63], Harray[45][63], Harray[46][63], Harray[47][63], Harray[48][63], Harray[49][63], Harray[50][63], Harray[51][63], Harray[52][63], Harray[53][63], Harray[54][63], Harray[55][63], Harray[56][63], Harray[57][63], Harray[58][63], Harray[59][63], Harray[60][63], Harray[61][63], Harray[62][63], Harray[63][63], Harray[64][63], Harray[65][63], Harray[66][63], Harray[67][63], Harray[68][63], Harray[69][63], Harray[70][63], Harray[71][63], Harray[72][63], Harray[73][63], Harray[74][63], Harray[75][63], Harray[76][63], Harray[77][63], Harray[78][63], Harray[79][63], Harray[80][63], Harray[81][63], Harray[82][63], Harray[83][63], Harray[84][63], Harray[85][63], Harray[86][63], Harray[87][63], Harray[88][63], Harray[89][63], Harray[90][63], Harray[91][63], Harray[92][63], Harray[93][63], Harray[94][63], Harray[95][63], Harray[96][63], Harray[97][63], Harray[98][63], Harray[99][63], Harray[100][63], Harray[101][63], Harray[102][63], Harray[103][63], Harray[104][63], Harray[105][63], Harray[106][63], Harray[107][63], Harray[108][63], Harray[109][63], Harray[110][63], Harray[111][63], Harray[112][63], Harray[113][63], Harray[114][63], Harray[115][63], Harray[116][63], Harray[117][63], Harray[118][63], Harray[119][63], Harray[120][63], Harray[121][63], Harray[122][63], Harray[123][63], Harray[124][63], Harray[125][63], Harray[126][63], Harray[127][63]};
assign h_col_64 = {Harray[0][64], Harray[1][64], Harray[2][64], Harray[3][64], Harray[4][64], Harray[5][64], Harray[6][64], Harray[7][64], Harray[8][64], Harray[9][64], Harray[10][64], Harray[11][64], Harray[12][64], Harray[13][64], Harray[14][64], Harray[15][64], Harray[16][64], Harray[17][64], Harray[18][64], Harray[19][64], Harray[20][64], Harray[21][64], Harray[22][64], Harray[23][64], Harray[24][64], Harray[25][64], Harray[26][64], Harray[27][64], Harray[28][64], Harray[29][64], Harray[30][64], Harray[31][64], Harray[32][64], Harray[33][64], Harray[34][64], Harray[35][64], Harray[36][64], Harray[37][64], Harray[38][64], Harray[39][64], Harray[40][64], Harray[41][64], Harray[42][64], Harray[43][64], Harray[44][64], Harray[45][64], Harray[46][64], Harray[47][64], Harray[48][64], Harray[49][64], Harray[50][64], Harray[51][64], Harray[52][64], Harray[53][64], Harray[54][64], Harray[55][64], Harray[56][64], Harray[57][64], Harray[58][64], Harray[59][64], Harray[60][64], Harray[61][64], Harray[62][64], Harray[63][64], Harray[64][64], Harray[65][64], Harray[66][64], Harray[67][64], Harray[68][64], Harray[69][64], Harray[70][64], Harray[71][64], Harray[72][64], Harray[73][64], Harray[74][64], Harray[75][64], Harray[76][64], Harray[77][64], Harray[78][64], Harray[79][64], Harray[80][64], Harray[81][64], Harray[82][64], Harray[83][64], Harray[84][64], Harray[85][64], Harray[86][64], Harray[87][64], Harray[88][64], Harray[89][64], Harray[90][64], Harray[91][64], Harray[92][64], Harray[93][64], Harray[94][64], Harray[95][64], Harray[96][64], Harray[97][64], Harray[98][64], Harray[99][64], Harray[100][64], Harray[101][64], Harray[102][64], Harray[103][64], Harray[104][64], Harray[105][64], Harray[106][64], Harray[107][64], Harray[108][64], Harray[109][64], Harray[110][64], Harray[111][64], Harray[112][64], Harray[113][64], Harray[114][64], Harray[115][64], Harray[116][64], Harray[117][64], Harray[118][64], Harray[119][64], Harray[120][64], Harray[121][64], Harray[122][64], Harray[123][64], Harray[124][64], Harray[125][64], Harray[126][64], Harray[127][64]};
assign h_col_65 = {Harray[0][65], Harray[1][65], Harray[2][65], Harray[3][65], Harray[4][65], Harray[5][65], Harray[6][65], Harray[7][65], Harray[8][65], Harray[9][65], Harray[10][65], Harray[11][65], Harray[12][65], Harray[13][65], Harray[14][65], Harray[15][65], Harray[16][65], Harray[17][65], Harray[18][65], Harray[19][65], Harray[20][65], Harray[21][65], Harray[22][65], Harray[23][65], Harray[24][65], Harray[25][65], Harray[26][65], Harray[27][65], Harray[28][65], Harray[29][65], Harray[30][65], Harray[31][65], Harray[32][65], Harray[33][65], Harray[34][65], Harray[35][65], Harray[36][65], Harray[37][65], Harray[38][65], Harray[39][65], Harray[40][65], Harray[41][65], Harray[42][65], Harray[43][65], Harray[44][65], Harray[45][65], Harray[46][65], Harray[47][65], Harray[48][65], Harray[49][65], Harray[50][65], Harray[51][65], Harray[52][65], Harray[53][65], Harray[54][65], Harray[55][65], Harray[56][65], Harray[57][65], Harray[58][65], Harray[59][65], Harray[60][65], Harray[61][65], Harray[62][65], Harray[63][65], Harray[64][65], Harray[65][65], Harray[66][65], Harray[67][65], Harray[68][65], Harray[69][65], Harray[70][65], Harray[71][65], Harray[72][65], Harray[73][65], Harray[74][65], Harray[75][65], Harray[76][65], Harray[77][65], Harray[78][65], Harray[79][65], Harray[80][65], Harray[81][65], Harray[82][65], Harray[83][65], Harray[84][65], Harray[85][65], Harray[86][65], Harray[87][65], Harray[88][65], Harray[89][65], Harray[90][65], Harray[91][65], Harray[92][65], Harray[93][65], Harray[94][65], Harray[95][65], Harray[96][65], Harray[97][65], Harray[98][65], Harray[99][65], Harray[100][65], Harray[101][65], Harray[102][65], Harray[103][65], Harray[104][65], Harray[105][65], Harray[106][65], Harray[107][65], Harray[108][65], Harray[109][65], Harray[110][65], Harray[111][65], Harray[112][65], Harray[113][65], Harray[114][65], Harray[115][65], Harray[116][65], Harray[117][65], Harray[118][65], Harray[119][65], Harray[120][65], Harray[121][65], Harray[122][65], Harray[123][65], Harray[124][65], Harray[125][65], Harray[126][65], Harray[127][65]};
assign h_col_66 = {Harray[0][66], Harray[1][66], Harray[2][66], Harray[3][66], Harray[4][66], Harray[5][66], Harray[6][66], Harray[7][66], Harray[8][66], Harray[9][66], Harray[10][66], Harray[11][66], Harray[12][66], Harray[13][66], Harray[14][66], Harray[15][66], Harray[16][66], Harray[17][66], Harray[18][66], Harray[19][66], Harray[20][66], Harray[21][66], Harray[22][66], Harray[23][66], Harray[24][66], Harray[25][66], Harray[26][66], Harray[27][66], Harray[28][66], Harray[29][66], Harray[30][66], Harray[31][66], Harray[32][66], Harray[33][66], Harray[34][66], Harray[35][66], Harray[36][66], Harray[37][66], Harray[38][66], Harray[39][66], Harray[40][66], Harray[41][66], Harray[42][66], Harray[43][66], Harray[44][66], Harray[45][66], Harray[46][66], Harray[47][66], Harray[48][66], Harray[49][66], Harray[50][66], Harray[51][66], Harray[52][66], Harray[53][66], Harray[54][66], Harray[55][66], Harray[56][66], Harray[57][66], Harray[58][66], Harray[59][66], Harray[60][66], Harray[61][66], Harray[62][66], Harray[63][66], Harray[64][66], Harray[65][66], Harray[66][66], Harray[67][66], Harray[68][66], Harray[69][66], Harray[70][66], Harray[71][66], Harray[72][66], Harray[73][66], Harray[74][66], Harray[75][66], Harray[76][66], Harray[77][66], Harray[78][66], Harray[79][66], Harray[80][66], Harray[81][66], Harray[82][66], Harray[83][66], Harray[84][66], Harray[85][66], Harray[86][66], Harray[87][66], Harray[88][66], Harray[89][66], Harray[90][66], Harray[91][66], Harray[92][66], Harray[93][66], Harray[94][66], Harray[95][66], Harray[96][66], Harray[97][66], Harray[98][66], Harray[99][66], Harray[100][66], Harray[101][66], Harray[102][66], Harray[103][66], Harray[104][66], Harray[105][66], Harray[106][66], Harray[107][66], Harray[108][66], Harray[109][66], Harray[110][66], Harray[111][66], Harray[112][66], Harray[113][66], Harray[114][66], Harray[115][66], Harray[116][66], Harray[117][66], Harray[118][66], Harray[119][66], Harray[120][66], Harray[121][66], Harray[122][66], Harray[123][66], Harray[124][66], Harray[125][66], Harray[126][66], Harray[127][66]};
assign h_col_67 = {Harray[0][67], Harray[1][67], Harray[2][67], Harray[3][67], Harray[4][67], Harray[5][67], Harray[6][67], Harray[7][67], Harray[8][67], Harray[9][67], Harray[10][67], Harray[11][67], Harray[12][67], Harray[13][67], Harray[14][67], Harray[15][67], Harray[16][67], Harray[17][67], Harray[18][67], Harray[19][67], Harray[20][67], Harray[21][67], Harray[22][67], Harray[23][67], Harray[24][67], Harray[25][67], Harray[26][67], Harray[27][67], Harray[28][67], Harray[29][67], Harray[30][67], Harray[31][67], Harray[32][67], Harray[33][67], Harray[34][67], Harray[35][67], Harray[36][67], Harray[37][67], Harray[38][67], Harray[39][67], Harray[40][67], Harray[41][67], Harray[42][67], Harray[43][67], Harray[44][67], Harray[45][67], Harray[46][67], Harray[47][67], Harray[48][67], Harray[49][67], Harray[50][67], Harray[51][67], Harray[52][67], Harray[53][67], Harray[54][67], Harray[55][67], Harray[56][67], Harray[57][67], Harray[58][67], Harray[59][67], Harray[60][67], Harray[61][67], Harray[62][67], Harray[63][67], Harray[64][67], Harray[65][67], Harray[66][67], Harray[67][67], Harray[68][67], Harray[69][67], Harray[70][67], Harray[71][67], Harray[72][67], Harray[73][67], Harray[74][67], Harray[75][67], Harray[76][67], Harray[77][67], Harray[78][67], Harray[79][67], Harray[80][67], Harray[81][67], Harray[82][67], Harray[83][67], Harray[84][67], Harray[85][67], Harray[86][67], Harray[87][67], Harray[88][67], Harray[89][67], Harray[90][67], Harray[91][67], Harray[92][67], Harray[93][67], Harray[94][67], Harray[95][67], Harray[96][67], Harray[97][67], Harray[98][67], Harray[99][67], Harray[100][67], Harray[101][67], Harray[102][67], Harray[103][67], Harray[104][67], Harray[105][67], Harray[106][67], Harray[107][67], Harray[108][67], Harray[109][67], Harray[110][67], Harray[111][67], Harray[112][67], Harray[113][67], Harray[114][67], Harray[115][67], Harray[116][67], Harray[117][67], Harray[118][67], Harray[119][67], Harray[120][67], Harray[121][67], Harray[122][67], Harray[123][67], Harray[124][67], Harray[125][67], Harray[126][67], Harray[127][67]};
assign h_col_68 = {Harray[0][68], Harray[1][68], Harray[2][68], Harray[3][68], Harray[4][68], Harray[5][68], Harray[6][68], Harray[7][68], Harray[8][68], Harray[9][68], Harray[10][68], Harray[11][68], Harray[12][68], Harray[13][68], Harray[14][68], Harray[15][68], Harray[16][68], Harray[17][68], Harray[18][68], Harray[19][68], Harray[20][68], Harray[21][68], Harray[22][68], Harray[23][68], Harray[24][68], Harray[25][68], Harray[26][68], Harray[27][68], Harray[28][68], Harray[29][68], Harray[30][68], Harray[31][68], Harray[32][68], Harray[33][68], Harray[34][68], Harray[35][68], Harray[36][68], Harray[37][68], Harray[38][68], Harray[39][68], Harray[40][68], Harray[41][68], Harray[42][68], Harray[43][68], Harray[44][68], Harray[45][68], Harray[46][68], Harray[47][68], Harray[48][68], Harray[49][68], Harray[50][68], Harray[51][68], Harray[52][68], Harray[53][68], Harray[54][68], Harray[55][68], Harray[56][68], Harray[57][68], Harray[58][68], Harray[59][68], Harray[60][68], Harray[61][68], Harray[62][68], Harray[63][68], Harray[64][68], Harray[65][68], Harray[66][68], Harray[67][68], Harray[68][68], Harray[69][68], Harray[70][68], Harray[71][68], Harray[72][68], Harray[73][68], Harray[74][68], Harray[75][68], Harray[76][68], Harray[77][68], Harray[78][68], Harray[79][68], Harray[80][68], Harray[81][68], Harray[82][68], Harray[83][68], Harray[84][68], Harray[85][68], Harray[86][68], Harray[87][68], Harray[88][68], Harray[89][68], Harray[90][68], Harray[91][68], Harray[92][68], Harray[93][68], Harray[94][68], Harray[95][68], Harray[96][68], Harray[97][68], Harray[98][68], Harray[99][68], Harray[100][68], Harray[101][68], Harray[102][68], Harray[103][68], Harray[104][68], Harray[105][68], Harray[106][68], Harray[107][68], Harray[108][68], Harray[109][68], Harray[110][68], Harray[111][68], Harray[112][68], Harray[113][68], Harray[114][68], Harray[115][68], Harray[116][68], Harray[117][68], Harray[118][68], Harray[119][68], Harray[120][68], Harray[121][68], Harray[122][68], Harray[123][68], Harray[124][68], Harray[125][68], Harray[126][68], Harray[127][68]};
assign h_col_69 = {Harray[0][69], Harray[1][69], Harray[2][69], Harray[3][69], Harray[4][69], Harray[5][69], Harray[6][69], Harray[7][69], Harray[8][69], Harray[9][69], Harray[10][69], Harray[11][69], Harray[12][69], Harray[13][69], Harray[14][69], Harray[15][69], Harray[16][69], Harray[17][69], Harray[18][69], Harray[19][69], Harray[20][69], Harray[21][69], Harray[22][69], Harray[23][69], Harray[24][69], Harray[25][69], Harray[26][69], Harray[27][69], Harray[28][69], Harray[29][69], Harray[30][69], Harray[31][69], Harray[32][69], Harray[33][69], Harray[34][69], Harray[35][69], Harray[36][69], Harray[37][69], Harray[38][69], Harray[39][69], Harray[40][69], Harray[41][69], Harray[42][69], Harray[43][69], Harray[44][69], Harray[45][69], Harray[46][69], Harray[47][69], Harray[48][69], Harray[49][69], Harray[50][69], Harray[51][69], Harray[52][69], Harray[53][69], Harray[54][69], Harray[55][69], Harray[56][69], Harray[57][69], Harray[58][69], Harray[59][69], Harray[60][69], Harray[61][69], Harray[62][69], Harray[63][69], Harray[64][69], Harray[65][69], Harray[66][69], Harray[67][69], Harray[68][69], Harray[69][69], Harray[70][69], Harray[71][69], Harray[72][69], Harray[73][69], Harray[74][69], Harray[75][69], Harray[76][69], Harray[77][69], Harray[78][69], Harray[79][69], Harray[80][69], Harray[81][69], Harray[82][69], Harray[83][69], Harray[84][69], Harray[85][69], Harray[86][69], Harray[87][69], Harray[88][69], Harray[89][69], Harray[90][69], Harray[91][69], Harray[92][69], Harray[93][69], Harray[94][69], Harray[95][69], Harray[96][69], Harray[97][69], Harray[98][69], Harray[99][69], Harray[100][69], Harray[101][69], Harray[102][69], Harray[103][69], Harray[104][69], Harray[105][69], Harray[106][69], Harray[107][69], Harray[108][69], Harray[109][69], Harray[110][69], Harray[111][69], Harray[112][69], Harray[113][69], Harray[114][69], Harray[115][69], Harray[116][69], Harray[117][69], Harray[118][69], Harray[119][69], Harray[120][69], Harray[121][69], Harray[122][69], Harray[123][69], Harray[124][69], Harray[125][69], Harray[126][69], Harray[127][69]};
assign h_col_70 = {Harray[0][70], Harray[1][70], Harray[2][70], Harray[3][70], Harray[4][70], Harray[5][70], Harray[6][70], Harray[7][70], Harray[8][70], Harray[9][70], Harray[10][70], Harray[11][70], Harray[12][70], Harray[13][70], Harray[14][70], Harray[15][70], Harray[16][70], Harray[17][70], Harray[18][70], Harray[19][70], Harray[20][70], Harray[21][70], Harray[22][70], Harray[23][70], Harray[24][70], Harray[25][70], Harray[26][70], Harray[27][70], Harray[28][70], Harray[29][70], Harray[30][70], Harray[31][70], Harray[32][70], Harray[33][70], Harray[34][70], Harray[35][70], Harray[36][70], Harray[37][70], Harray[38][70], Harray[39][70], Harray[40][70], Harray[41][70], Harray[42][70], Harray[43][70], Harray[44][70], Harray[45][70], Harray[46][70], Harray[47][70], Harray[48][70], Harray[49][70], Harray[50][70], Harray[51][70], Harray[52][70], Harray[53][70], Harray[54][70], Harray[55][70], Harray[56][70], Harray[57][70], Harray[58][70], Harray[59][70], Harray[60][70], Harray[61][70], Harray[62][70], Harray[63][70], Harray[64][70], Harray[65][70], Harray[66][70], Harray[67][70], Harray[68][70], Harray[69][70], Harray[70][70], Harray[71][70], Harray[72][70], Harray[73][70], Harray[74][70], Harray[75][70], Harray[76][70], Harray[77][70], Harray[78][70], Harray[79][70], Harray[80][70], Harray[81][70], Harray[82][70], Harray[83][70], Harray[84][70], Harray[85][70], Harray[86][70], Harray[87][70], Harray[88][70], Harray[89][70], Harray[90][70], Harray[91][70], Harray[92][70], Harray[93][70], Harray[94][70], Harray[95][70], Harray[96][70], Harray[97][70], Harray[98][70], Harray[99][70], Harray[100][70], Harray[101][70], Harray[102][70], Harray[103][70], Harray[104][70], Harray[105][70], Harray[106][70], Harray[107][70], Harray[108][70], Harray[109][70], Harray[110][70], Harray[111][70], Harray[112][70], Harray[113][70], Harray[114][70], Harray[115][70], Harray[116][70], Harray[117][70], Harray[118][70], Harray[119][70], Harray[120][70], Harray[121][70], Harray[122][70], Harray[123][70], Harray[124][70], Harray[125][70], Harray[126][70], Harray[127][70]};
assign h_col_71 = {Harray[0][71], Harray[1][71], Harray[2][71], Harray[3][71], Harray[4][71], Harray[5][71], Harray[6][71], Harray[7][71], Harray[8][71], Harray[9][71], Harray[10][71], Harray[11][71], Harray[12][71], Harray[13][71], Harray[14][71], Harray[15][71], Harray[16][71], Harray[17][71], Harray[18][71], Harray[19][71], Harray[20][71], Harray[21][71], Harray[22][71], Harray[23][71], Harray[24][71], Harray[25][71], Harray[26][71], Harray[27][71], Harray[28][71], Harray[29][71], Harray[30][71], Harray[31][71], Harray[32][71], Harray[33][71], Harray[34][71], Harray[35][71], Harray[36][71], Harray[37][71], Harray[38][71], Harray[39][71], Harray[40][71], Harray[41][71], Harray[42][71], Harray[43][71], Harray[44][71], Harray[45][71], Harray[46][71], Harray[47][71], Harray[48][71], Harray[49][71], Harray[50][71], Harray[51][71], Harray[52][71], Harray[53][71], Harray[54][71], Harray[55][71], Harray[56][71], Harray[57][71], Harray[58][71], Harray[59][71], Harray[60][71], Harray[61][71], Harray[62][71], Harray[63][71], Harray[64][71], Harray[65][71], Harray[66][71], Harray[67][71], Harray[68][71], Harray[69][71], Harray[70][71], Harray[71][71], Harray[72][71], Harray[73][71], Harray[74][71], Harray[75][71], Harray[76][71], Harray[77][71], Harray[78][71], Harray[79][71], Harray[80][71], Harray[81][71], Harray[82][71], Harray[83][71], Harray[84][71], Harray[85][71], Harray[86][71], Harray[87][71], Harray[88][71], Harray[89][71], Harray[90][71], Harray[91][71], Harray[92][71], Harray[93][71], Harray[94][71], Harray[95][71], Harray[96][71], Harray[97][71], Harray[98][71], Harray[99][71], Harray[100][71], Harray[101][71], Harray[102][71], Harray[103][71], Harray[104][71], Harray[105][71], Harray[106][71], Harray[107][71], Harray[108][71], Harray[109][71], Harray[110][71], Harray[111][71], Harray[112][71], Harray[113][71], Harray[114][71], Harray[115][71], Harray[116][71], Harray[117][71], Harray[118][71], Harray[119][71], Harray[120][71], Harray[121][71], Harray[122][71], Harray[123][71], Harray[124][71], Harray[125][71], Harray[126][71], Harray[127][71]};
assign h_col_72 = {Harray[0][72], Harray[1][72], Harray[2][72], Harray[3][72], Harray[4][72], Harray[5][72], Harray[6][72], Harray[7][72], Harray[8][72], Harray[9][72], Harray[10][72], Harray[11][72], Harray[12][72], Harray[13][72], Harray[14][72], Harray[15][72], Harray[16][72], Harray[17][72], Harray[18][72], Harray[19][72], Harray[20][72], Harray[21][72], Harray[22][72], Harray[23][72], Harray[24][72], Harray[25][72], Harray[26][72], Harray[27][72], Harray[28][72], Harray[29][72], Harray[30][72], Harray[31][72], Harray[32][72], Harray[33][72], Harray[34][72], Harray[35][72], Harray[36][72], Harray[37][72], Harray[38][72], Harray[39][72], Harray[40][72], Harray[41][72], Harray[42][72], Harray[43][72], Harray[44][72], Harray[45][72], Harray[46][72], Harray[47][72], Harray[48][72], Harray[49][72], Harray[50][72], Harray[51][72], Harray[52][72], Harray[53][72], Harray[54][72], Harray[55][72], Harray[56][72], Harray[57][72], Harray[58][72], Harray[59][72], Harray[60][72], Harray[61][72], Harray[62][72], Harray[63][72], Harray[64][72], Harray[65][72], Harray[66][72], Harray[67][72], Harray[68][72], Harray[69][72], Harray[70][72], Harray[71][72], Harray[72][72], Harray[73][72], Harray[74][72], Harray[75][72], Harray[76][72], Harray[77][72], Harray[78][72], Harray[79][72], Harray[80][72], Harray[81][72], Harray[82][72], Harray[83][72], Harray[84][72], Harray[85][72], Harray[86][72], Harray[87][72], Harray[88][72], Harray[89][72], Harray[90][72], Harray[91][72], Harray[92][72], Harray[93][72], Harray[94][72], Harray[95][72], Harray[96][72], Harray[97][72], Harray[98][72], Harray[99][72], Harray[100][72], Harray[101][72], Harray[102][72], Harray[103][72], Harray[104][72], Harray[105][72], Harray[106][72], Harray[107][72], Harray[108][72], Harray[109][72], Harray[110][72], Harray[111][72], Harray[112][72], Harray[113][72], Harray[114][72], Harray[115][72], Harray[116][72], Harray[117][72], Harray[118][72], Harray[119][72], Harray[120][72], Harray[121][72], Harray[122][72], Harray[123][72], Harray[124][72], Harray[125][72], Harray[126][72], Harray[127][72]};
assign h_col_73 = {Harray[0][73], Harray[1][73], Harray[2][73], Harray[3][73], Harray[4][73], Harray[5][73], Harray[6][73], Harray[7][73], Harray[8][73], Harray[9][73], Harray[10][73], Harray[11][73], Harray[12][73], Harray[13][73], Harray[14][73], Harray[15][73], Harray[16][73], Harray[17][73], Harray[18][73], Harray[19][73], Harray[20][73], Harray[21][73], Harray[22][73], Harray[23][73], Harray[24][73], Harray[25][73], Harray[26][73], Harray[27][73], Harray[28][73], Harray[29][73], Harray[30][73], Harray[31][73], Harray[32][73], Harray[33][73], Harray[34][73], Harray[35][73], Harray[36][73], Harray[37][73], Harray[38][73], Harray[39][73], Harray[40][73], Harray[41][73], Harray[42][73], Harray[43][73], Harray[44][73], Harray[45][73], Harray[46][73], Harray[47][73], Harray[48][73], Harray[49][73], Harray[50][73], Harray[51][73], Harray[52][73], Harray[53][73], Harray[54][73], Harray[55][73], Harray[56][73], Harray[57][73], Harray[58][73], Harray[59][73], Harray[60][73], Harray[61][73], Harray[62][73], Harray[63][73], Harray[64][73], Harray[65][73], Harray[66][73], Harray[67][73], Harray[68][73], Harray[69][73], Harray[70][73], Harray[71][73], Harray[72][73], Harray[73][73], Harray[74][73], Harray[75][73], Harray[76][73], Harray[77][73], Harray[78][73], Harray[79][73], Harray[80][73], Harray[81][73], Harray[82][73], Harray[83][73], Harray[84][73], Harray[85][73], Harray[86][73], Harray[87][73], Harray[88][73], Harray[89][73], Harray[90][73], Harray[91][73], Harray[92][73], Harray[93][73], Harray[94][73], Harray[95][73], Harray[96][73], Harray[97][73], Harray[98][73], Harray[99][73], Harray[100][73], Harray[101][73], Harray[102][73], Harray[103][73], Harray[104][73], Harray[105][73], Harray[106][73], Harray[107][73], Harray[108][73], Harray[109][73], Harray[110][73], Harray[111][73], Harray[112][73], Harray[113][73], Harray[114][73], Harray[115][73], Harray[116][73], Harray[117][73], Harray[118][73], Harray[119][73], Harray[120][73], Harray[121][73], Harray[122][73], Harray[123][73], Harray[124][73], Harray[125][73], Harray[126][73], Harray[127][73]};
assign h_col_74 = {Harray[0][74], Harray[1][74], Harray[2][74], Harray[3][74], Harray[4][74], Harray[5][74], Harray[6][74], Harray[7][74], Harray[8][74], Harray[9][74], Harray[10][74], Harray[11][74], Harray[12][74], Harray[13][74], Harray[14][74], Harray[15][74], Harray[16][74], Harray[17][74], Harray[18][74], Harray[19][74], Harray[20][74], Harray[21][74], Harray[22][74], Harray[23][74], Harray[24][74], Harray[25][74], Harray[26][74], Harray[27][74], Harray[28][74], Harray[29][74], Harray[30][74], Harray[31][74], Harray[32][74], Harray[33][74], Harray[34][74], Harray[35][74], Harray[36][74], Harray[37][74], Harray[38][74], Harray[39][74], Harray[40][74], Harray[41][74], Harray[42][74], Harray[43][74], Harray[44][74], Harray[45][74], Harray[46][74], Harray[47][74], Harray[48][74], Harray[49][74], Harray[50][74], Harray[51][74], Harray[52][74], Harray[53][74], Harray[54][74], Harray[55][74], Harray[56][74], Harray[57][74], Harray[58][74], Harray[59][74], Harray[60][74], Harray[61][74], Harray[62][74], Harray[63][74], Harray[64][74], Harray[65][74], Harray[66][74], Harray[67][74], Harray[68][74], Harray[69][74], Harray[70][74], Harray[71][74], Harray[72][74], Harray[73][74], Harray[74][74], Harray[75][74], Harray[76][74], Harray[77][74], Harray[78][74], Harray[79][74], Harray[80][74], Harray[81][74], Harray[82][74], Harray[83][74], Harray[84][74], Harray[85][74], Harray[86][74], Harray[87][74], Harray[88][74], Harray[89][74], Harray[90][74], Harray[91][74], Harray[92][74], Harray[93][74], Harray[94][74], Harray[95][74], Harray[96][74], Harray[97][74], Harray[98][74], Harray[99][74], Harray[100][74], Harray[101][74], Harray[102][74], Harray[103][74], Harray[104][74], Harray[105][74], Harray[106][74], Harray[107][74], Harray[108][74], Harray[109][74], Harray[110][74], Harray[111][74], Harray[112][74], Harray[113][74], Harray[114][74], Harray[115][74], Harray[116][74], Harray[117][74], Harray[118][74], Harray[119][74], Harray[120][74], Harray[121][74], Harray[122][74], Harray[123][74], Harray[124][74], Harray[125][74], Harray[126][74], Harray[127][74]};
assign h_col_75 = {Harray[0][75], Harray[1][75], Harray[2][75], Harray[3][75], Harray[4][75], Harray[5][75], Harray[6][75], Harray[7][75], Harray[8][75], Harray[9][75], Harray[10][75], Harray[11][75], Harray[12][75], Harray[13][75], Harray[14][75], Harray[15][75], Harray[16][75], Harray[17][75], Harray[18][75], Harray[19][75], Harray[20][75], Harray[21][75], Harray[22][75], Harray[23][75], Harray[24][75], Harray[25][75], Harray[26][75], Harray[27][75], Harray[28][75], Harray[29][75], Harray[30][75], Harray[31][75], Harray[32][75], Harray[33][75], Harray[34][75], Harray[35][75], Harray[36][75], Harray[37][75], Harray[38][75], Harray[39][75], Harray[40][75], Harray[41][75], Harray[42][75], Harray[43][75], Harray[44][75], Harray[45][75], Harray[46][75], Harray[47][75], Harray[48][75], Harray[49][75], Harray[50][75], Harray[51][75], Harray[52][75], Harray[53][75], Harray[54][75], Harray[55][75], Harray[56][75], Harray[57][75], Harray[58][75], Harray[59][75], Harray[60][75], Harray[61][75], Harray[62][75], Harray[63][75], Harray[64][75], Harray[65][75], Harray[66][75], Harray[67][75], Harray[68][75], Harray[69][75], Harray[70][75], Harray[71][75], Harray[72][75], Harray[73][75], Harray[74][75], Harray[75][75], Harray[76][75], Harray[77][75], Harray[78][75], Harray[79][75], Harray[80][75], Harray[81][75], Harray[82][75], Harray[83][75], Harray[84][75], Harray[85][75], Harray[86][75], Harray[87][75], Harray[88][75], Harray[89][75], Harray[90][75], Harray[91][75], Harray[92][75], Harray[93][75], Harray[94][75], Harray[95][75], Harray[96][75], Harray[97][75], Harray[98][75], Harray[99][75], Harray[100][75], Harray[101][75], Harray[102][75], Harray[103][75], Harray[104][75], Harray[105][75], Harray[106][75], Harray[107][75], Harray[108][75], Harray[109][75], Harray[110][75], Harray[111][75], Harray[112][75], Harray[113][75], Harray[114][75], Harray[115][75], Harray[116][75], Harray[117][75], Harray[118][75], Harray[119][75], Harray[120][75], Harray[121][75], Harray[122][75], Harray[123][75], Harray[124][75], Harray[125][75], Harray[126][75], Harray[127][75]};
assign h_col_76 = {Harray[0][76], Harray[1][76], Harray[2][76], Harray[3][76], Harray[4][76], Harray[5][76], Harray[6][76], Harray[7][76], Harray[8][76], Harray[9][76], Harray[10][76], Harray[11][76], Harray[12][76], Harray[13][76], Harray[14][76], Harray[15][76], Harray[16][76], Harray[17][76], Harray[18][76], Harray[19][76], Harray[20][76], Harray[21][76], Harray[22][76], Harray[23][76], Harray[24][76], Harray[25][76], Harray[26][76], Harray[27][76], Harray[28][76], Harray[29][76], Harray[30][76], Harray[31][76], Harray[32][76], Harray[33][76], Harray[34][76], Harray[35][76], Harray[36][76], Harray[37][76], Harray[38][76], Harray[39][76], Harray[40][76], Harray[41][76], Harray[42][76], Harray[43][76], Harray[44][76], Harray[45][76], Harray[46][76], Harray[47][76], Harray[48][76], Harray[49][76], Harray[50][76], Harray[51][76], Harray[52][76], Harray[53][76], Harray[54][76], Harray[55][76], Harray[56][76], Harray[57][76], Harray[58][76], Harray[59][76], Harray[60][76], Harray[61][76], Harray[62][76], Harray[63][76], Harray[64][76], Harray[65][76], Harray[66][76], Harray[67][76], Harray[68][76], Harray[69][76], Harray[70][76], Harray[71][76], Harray[72][76], Harray[73][76], Harray[74][76], Harray[75][76], Harray[76][76], Harray[77][76], Harray[78][76], Harray[79][76], Harray[80][76], Harray[81][76], Harray[82][76], Harray[83][76], Harray[84][76], Harray[85][76], Harray[86][76], Harray[87][76], Harray[88][76], Harray[89][76], Harray[90][76], Harray[91][76], Harray[92][76], Harray[93][76], Harray[94][76], Harray[95][76], Harray[96][76], Harray[97][76], Harray[98][76], Harray[99][76], Harray[100][76], Harray[101][76], Harray[102][76], Harray[103][76], Harray[104][76], Harray[105][76], Harray[106][76], Harray[107][76], Harray[108][76], Harray[109][76], Harray[110][76], Harray[111][76], Harray[112][76], Harray[113][76], Harray[114][76], Harray[115][76], Harray[116][76], Harray[117][76], Harray[118][76], Harray[119][76], Harray[120][76], Harray[121][76], Harray[122][76], Harray[123][76], Harray[124][76], Harray[125][76], Harray[126][76], Harray[127][76]};
assign h_col_77 = {Harray[0][77], Harray[1][77], Harray[2][77], Harray[3][77], Harray[4][77], Harray[5][77], Harray[6][77], Harray[7][77], Harray[8][77], Harray[9][77], Harray[10][77], Harray[11][77], Harray[12][77], Harray[13][77], Harray[14][77], Harray[15][77], Harray[16][77], Harray[17][77], Harray[18][77], Harray[19][77], Harray[20][77], Harray[21][77], Harray[22][77], Harray[23][77], Harray[24][77], Harray[25][77], Harray[26][77], Harray[27][77], Harray[28][77], Harray[29][77], Harray[30][77], Harray[31][77], Harray[32][77], Harray[33][77], Harray[34][77], Harray[35][77], Harray[36][77], Harray[37][77], Harray[38][77], Harray[39][77], Harray[40][77], Harray[41][77], Harray[42][77], Harray[43][77], Harray[44][77], Harray[45][77], Harray[46][77], Harray[47][77], Harray[48][77], Harray[49][77], Harray[50][77], Harray[51][77], Harray[52][77], Harray[53][77], Harray[54][77], Harray[55][77], Harray[56][77], Harray[57][77], Harray[58][77], Harray[59][77], Harray[60][77], Harray[61][77], Harray[62][77], Harray[63][77], Harray[64][77], Harray[65][77], Harray[66][77], Harray[67][77], Harray[68][77], Harray[69][77], Harray[70][77], Harray[71][77], Harray[72][77], Harray[73][77], Harray[74][77], Harray[75][77], Harray[76][77], Harray[77][77], Harray[78][77], Harray[79][77], Harray[80][77], Harray[81][77], Harray[82][77], Harray[83][77], Harray[84][77], Harray[85][77], Harray[86][77], Harray[87][77], Harray[88][77], Harray[89][77], Harray[90][77], Harray[91][77], Harray[92][77], Harray[93][77], Harray[94][77], Harray[95][77], Harray[96][77], Harray[97][77], Harray[98][77], Harray[99][77], Harray[100][77], Harray[101][77], Harray[102][77], Harray[103][77], Harray[104][77], Harray[105][77], Harray[106][77], Harray[107][77], Harray[108][77], Harray[109][77], Harray[110][77], Harray[111][77], Harray[112][77], Harray[113][77], Harray[114][77], Harray[115][77], Harray[116][77], Harray[117][77], Harray[118][77], Harray[119][77], Harray[120][77], Harray[121][77], Harray[122][77], Harray[123][77], Harray[124][77], Harray[125][77], Harray[126][77], Harray[127][77]};
assign h_col_78 = {Harray[0][78], Harray[1][78], Harray[2][78], Harray[3][78], Harray[4][78], Harray[5][78], Harray[6][78], Harray[7][78], Harray[8][78], Harray[9][78], Harray[10][78], Harray[11][78], Harray[12][78], Harray[13][78], Harray[14][78], Harray[15][78], Harray[16][78], Harray[17][78], Harray[18][78], Harray[19][78], Harray[20][78], Harray[21][78], Harray[22][78], Harray[23][78], Harray[24][78], Harray[25][78], Harray[26][78], Harray[27][78], Harray[28][78], Harray[29][78], Harray[30][78], Harray[31][78], Harray[32][78], Harray[33][78], Harray[34][78], Harray[35][78], Harray[36][78], Harray[37][78], Harray[38][78], Harray[39][78], Harray[40][78], Harray[41][78], Harray[42][78], Harray[43][78], Harray[44][78], Harray[45][78], Harray[46][78], Harray[47][78], Harray[48][78], Harray[49][78], Harray[50][78], Harray[51][78], Harray[52][78], Harray[53][78], Harray[54][78], Harray[55][78], Harray[56][78], Harray[57][78], Harray[58][78], Harray[59][78], Harray[60][78], Harray[61][78], Harray[62][78], Harray[63][78], Harray[64][78], Harray[65][78], Harray[66][78], Harray[67][78], Harray[68][78], Harray[69][78], Harray[70][78], Harray[71][78], Harray[72][78], Harray[73][78], Harray[74][78], Harray[75][78], Harray[76][78], Harray[77][78], Harray[78][78], Harray[79][78], Harray[80][78], Harray[81][78], Harray[82][78], Harray[83][78], Harray[84][78], Harray[85][78], Harray[86][78], Harray[87][78], Harray[88][78], Harray[89][78], Harray[90][78], Harray[91][78], Harray[92][78], Harray[93][78], Harray[94][78], Harray[95][78], Harray[96][78], Harray[97][78], Harray[98][78], Harray[99][78], Harray[100][78], Harray[101][78], Harray[102][78], Harray[103][78], Harray[104][78], Harray[105][78], Harray[106][78], Harray[107][78], Harray[108][78], Harray[109][78], Harray[110][78], Harray[111][78], Harray[112][78], Harray[113][78], Harray[114][78], Harray[115][78], Harray[116][78], Harray[117][78], Harray[118][78], Harray[119][78], Harray[120][78], Harray[121][78], Harray[122][78], Harray[123][78], Harray[124][78], Harray[125][78], Harray[126][78], Harray[127][78]};
assign h_col_79 = {Harray[0][79], Harray[1][79], Harray[2][79], Harray[3][79], Harray[4][79], Harray[5][79], Harray[6][79], Harray[7][79], Harray[8][79], Harray[9][79], Harray[10][79], Harray[11][79], Harray[12][79], Harray[13][79], Harray[14][79], Harray[15][79], Harray[16][79], Harray[17][79], Harray[18][79], Harray[19][79], Harray[20][79], Harray[21][79], Harray[22][79], Harray[23][79], Harray[24][79], Harray[25][79], Harray[26][79], Harray[27][79], Harray[28][79], Harray[29][79], Harray[30][79], Harray[31][79], Harray[32][79], Harray[33][79], Harray[34][79], Harray[35][79], Harray[36][79], Harray[37][79], Harray[38][79], Harray[39][79], Harray[40][79], Harray[41][79], Harray[42][79], Harray[43][79], Harray[44][79], Harray[45][79], Harray[46][79], Harray[47][79], Harray[48][79], Harray[49][79], Harray[50][79], Harray[51][79], Harray[52][79], Harray[53][79], Harray[54][79], Harray[55][79], Harray[56][79], Harray[57][79], Harray[58][79], Harray[59][79], Harray[60][79], Harray[61][79], Harray[62][79], Harray[63][79], Harray[64][79], Harray[65][79], Harray[66][79], Harray[67][79], Harray[68][79], Harray[69][79], Harray[70][79], Harray[71][79], Harray[72][79], Harray[73][79], Harray[74][79], Harray[75][79], Harray[76][79], Harray[77][79], Harray[78][79], Harray[79][79], Harray[80][79], Harray[81][79], Harray[82][79], Harray[83][79], Harray[84][79], Harray[85][79], Harray[86][79], Harray[87][79], Harray[88][79], Harray[89][79], Harray[90][79], Harray[91][79], Harray[92][79], Harray[93][79], Harray[94][79], Harray[95][79], Harray[96][79], Harray[97][79], Harray[98][79], Harray[99][79], Harray[100][79], Harray[101][79], Harray[102][79], Harray[103][79], Harray[104][79], Harray[105][79], Harray[106][79], Harray[107][79], Harray[108][79], Harray[109][79], Harray[110][79], Harray[111][79], Harray[112][79], Harray[113][79], Harray[114][79], Harray[115][79], Harray[116][79], Harray[117][79], Harray[118][79], Harray[119][79], Harray[120][79], Harray[121][79], Harray[122][79], Harray[123][79], Harray[124][79], Harray[125][79], Harray[126][79], Harray[127][79]};
assign h_col_80 = {Harray[0][80], Harray[1][80], Harray[2][80], Harray[3][80], Harray[4][80], Harray[5][80], Harray[6][80], Harray[7][80], Harray[8][80], Harray[9][80], Harray[10][80], Harray[11][80], Harray[12][80], Harray[13][80], Harray[14][80], Harray[15][80], Harray[16][80], Harray[17][80], Harray[18][80], Harray[19][80], Harray[20][80], Harray[21][80], Harray[22][80], Harray[23][80], Harray[24][80], Harray[25][80], Harray[26][80], Harray[27][80], Harray[28][80], Harray[29][80], Harray[30][80], Harray[31][80], Harray[32][80], Harray[33][80], Harray[34][80], Harray[35][80], Harray[36][80], Harray[37][80], Harray[38][80], Harray[39][80], Harray[40][80], Harray[41][80], Harray[42][80], Harray[43][80], Harray[44][80], Harray[45][80], Harray[46][80], Harray[47][80], Harray[48][80], Harray[49][80], Harray[50][80], Harray[51][80], Harray[52][80], Harray[53][80], Harray[54][80], Harray[55][80], Harray[56][80], Harray[57][80], Harray[58][80], Harray[59][80], Harray[60][80], Harray[61][80], Harray[62][80], Harray[63][80], Harray[64][80], Harray[65][80], Harray[66][80], Harray[67][80], Harray[68][80], Harray[69][80], Harray[70][80], Harray[71][80], Harray[72][80], Harray[73][80], Harray[74][80], Harray[75][80], Harray[76][80], Harray[77][80], Harray[78][80], Harray[79][80], Harray[80][80], Harray[81][80], Harray[82][80], Harray[83][80], Harray[84][80], Harray[85][80], Harray[86][80], Harray[87][80], Harray[88][80], Harray[89][80], Harray[90][80], Harray[91][80], Harray[92][80], Harray[93][80], Harray[94][80], Harray[95][80], Harray[96][80], Harray[97][80], Harray[98][80], Harray[99][80], Harray[100][80], Harray[101][80], Harray[102][80], Harray[103][80], Harray[104][80], Harray[105][80], Harray[106][80], Harray[107][80], Harray[108][80], Harray[109][80], Harray[110][80], Harray[111][80], Harray[112][80], Harray[113][80], Harray[114][80], Harray[115][80], Harray[116][80], Harray[117][80], Harray[118][80], Harray[119][80], Harray[120][80], Harray[121][80], Harray[122][80], Harray[123][80], Harray[124][80], Harray[125][80], Harray[126][80], Harray[127][80]};
assign h_col_81 = {Harray[0][81], Harray[1][81], Harray[2][81], Harray[3][81], Harray[4][81], Harray[5][81], Harray[6][81], Harray[7][81], Harray[8][81], Harray[9][81], Harray[10][81], Harray[11][81], Harray[12][81], Harray[13][81], Harray[14][81], Harray[15][81], Harray[16][81], Harray[17][81], Harray[18][81], Harray[19][81], Harray[20][81], Harray[21][81], Harray[22][81], Harray[23][81], Harray[24][81], Harray[25][81], Harray[26][81], Harray[27][81], Harray[28][81], Harray[29][81], Harray[30][81], Harray[31][81], Harray[32][81], Harray[33][81], Harray[34][81], Harray[35][81], Harray[36][81], Harray[37][81], Harray[38][81], Harray[39][81], Harray[40][81], Harray[41][81], Harray[42][81], Harray[43][81], Harray[44][81], Harray[45][81], Harray[46][81], Harray[47][81], Harray[48][81], Harray[49][81], Harray[50][81], Harray[51][81], Harray[52][81], Harray[53][81], Harray[54][81], Harray[55][81], Harray[56][81], Harray[57][81], Harray[58][81], Harray[59][81], Harray[60][81], Harray[61][81], Harray[62][81], Harray[63][81], Harray[64][81], Harray[65][81], Harray[66][81], Harray[67][81], Harray[68][81], Harray[69][81], Harray[70][81], Harray[71][81], Harray[72][81], Harray[73][81], Harray[74][81], Harray[75][81], Harray[76][81], Harray[77][81], Harray[78][81], Harray[79][81], Harray[80][81], Harray[81][81], Harray[82][81], Harray[83][81], Harray[84][81], Harray[85][81], Harray[86][81], Harray[87][81], Harray[88][81], Harray[89][81], Harray[90][81], Harray[91][81], Harray[92][81], Harray[93][81], Harray[94][81], Harray[95][81], Harray[96][81], Harray[97][81], Harray[98][81], Harray[99][81], Harray[100][81], Harray[101][81], Harray[102][81], Harray[103][81], Harray[104][81], Harray[105][81], Harray[106][81], Harray[107][81], Harray[108][81], Harray[109][81], Harray[110][81], Harray[111][81], Harray[112][81], Harray[113][81], Harray[114][81], Harray[115][81], Harray[116][81], Harray[117][81], Harray[118][81], Harray[119][81], Harray[120][81], Harray[121][81], Harray[122][81], Harray[123][81], Harray[124][81], Harray[125][81], Harray[126][81], Harray[127][81]};
assign h_col_82 = {Harray[0][82], Harray[1][82], Harray[2][82], Harray[3][82], Harray[4][82], Harray[5][82], Harray[6][82], Harray[7][82], Harray[8][82], Harray[9][82], Harray[10][82], Harray[11][82], Harray[12][82], Harray[13][82], Harray[14][82], Harray[15][82], Harray[16][82], Harray[17][82], Harray[18][82], Harray[19][82], Harray[20][82], Harray[21][82], Harray[22][82], Harray[23][82], Harray[24][82], Harray[25][82], Harray[26][82], Harray[27][82], Harray[28][82], Harray[29][82], Harray[30][82], Harray[31][82], Harray[32][82], Harray[33][82], Harray[34][82], Harray[35][82], Harray[36][82], Harray[37][82], Harray[38][82], Harray[39][82], Harray[40][82], Harray[41][82], Harray[42][82], Harray[43][82], Harray[44][82], Harray[45][82], Harray[46][82], Harray[47][82], Harray[48][82], Harray[49][82], Harray[50][82], Harray[51][82], Harray[52][82], Harray[53][82], Harray[54][82], Harray[55][82], Harray[56][82], Harray[57][82], Harray[58][82], Harray[59][82], Harray[60][82], Harray[61][82], Harray[62][82], Harray[63][82], Harray[64][82], Harray[65][82], Harray[66][82], Harray[67][82], Harray[68][82], Harray[69][82], Harray[70][82], Harray[71][82], Harray[72][82], Harray[73][82], Harray[74][82], Harray[75][82], Harray[76][82], Harray[77][82], Harray[78][82], Harray[79][82], Harray[80][82], Harray[81][82], Harray[82][82], Harray[83][82], Harray[84][82], Harray[85][82], Harray[86][82], Harray[87][82], Harray[88][82], Harray[89][82], Harray[90][82], Harray[91][82], Harray[92][82], Harray[93][82], Harray[94][82], Harray[95][82], Harray[96][82], Harray[97][82], Harray[98][82], Harray[99][82], Harray[100][82], Harray[101][82], Harray[102][82], Harray[103][82], Harray[104][82], Harray[105][82], Harray[106][82], Harray[107][82], Harray[108][82], Harray[109][82], Harray[110][82], Harray[111][82], Harray[112][82], Harray[113][82], Harray[114][82], Harray[115][82], Harray[116][82], Harray[117][82], Harray[118][82], Harray[119][82], Harray[120][82], Harray[121][82], Harray[122][82], Harray[123][82], Harray[124][82], Harray[125][82], Harray[126][82], Harray[127][82]};
assign h_col_83 = {Harray[0][83], Harray[1][83], Harray[2][83], Harray[3][83], Harray[4][83], Harray[5][83], Harray[6][83], Harray[7][83], Harray[8][83], Harray[9][83], Harray[10][83], Harray[11][83], Harray[12][83], Harray[13][83], Harray[14][83], Harray[15][83], Harray[16][83], Harray[17][83], Harray[18][83], Harray[19][83], Harray[20][83], Harray[21][83], Harray[22][83], Harray[23][83], Harray[24][83], Harray[25][83], Harray[26][83], Harray[27][83], Harray[28][83], Harray[29][83], Harray[30][83], Harray[31][83], Harray[32][83], Harray[33][83], Harray[34][83], Harray[35][83], Harray[36][83], Harray[37][83], Harray[38][83], Harray[39][83], Harray[40][83], Harray[41][83], Harray[42][83], Harray[43][83], Harray[44][83], Harray[45][83], Harray[46][83], Harray[47][83], Harray[48][83], Harray[49][83], Harray[50][83], Harray[51][83], Harray[52][83], Harray[53][83], Harray[54][83], Harray[55][83], Harray[56][83], Harray[57][83], Harray[58][83], Harray[59][83], Harray[60][83], Harray[61][83], Harray[62][83], Harray[63][83], Harray[64][83], Harray[65][83], Harray[66][83], Harray[67][83], Harray[68][83], Harray[69][83], Harray[70][83], Harray[71][83], Harray[72][83], Harray[73][83], Harray[74][83], Harray[75][83], Harray[76][83], Harray[77][83], Harray[78][83], Harray[79][83], Harray[80][83], Harray[81][83], Harray[82][83], Harray[83][83], Harray[84][83], Harray[85][83], Harray[86][83], Harray[87][83], Harray[88][83], Harray[89][83], Harray[90][83], Harray[91][83], Harray[92][83], Harray[93][83], Harray[94][83], Harray[95][83], Harray[96][83], Harray[97][83], Harray[98][83], Harray[99][83], Harray[100][83], Harray[101][83], Harray[102][83], Harray[103][83], Harray[104][83], Harray[105][83], Harray[106][83], Harray[107][83], Harray[108][83], Harray[109][83], Harray[110][83], Harray[111][83], Harray[112][83], Harray[113][83], Harray[114][83], Harray[115][83], Harray[116][83], Harray[117][83], Harray[118][83], Harray[119][83], Harray[120][83], Harray[121][83], Harray[122][83], Harray[123][83], Harray[124][83], Harray[125][83], Harray[126][83], Harray[127][83]};
assign h_col_84 = {Harray[0][84], Harray[1][84], Harray[2][84], Harray[3][84], Harray[4][84], Harray[5][84], Harray[6][84], Harray[7][84], Harray[8][84], Harray[9][84], Harray[10][84], Harray[11][84], Harray[12][84], Harray[13][84], Harray[14][84], Harray[15][84], Harray[16][84], Harray[17][84], Harray[18][84], Harray[19][84], Harray[20][84], Harray[21][84], Harray[22][84], Harray[23][84], Harray[24][84], Harray[25][84], Harray[26][84], Harray[27][84], Harray[28][84], Harray[29][84], Harray[30][84], Harray[31][84], Harray[32][84], Harray[33][84], Harray[34][84], Harray[35][84], Harray[36][84], Harray[37][84], Harray[38][84], Harray[39][84], Harray[40][84], Harray[41][84], Harray[42][84], Harray[43][84], Harray[44][84], Harray[45][84], Harray[46][84], Harray[47][84], Harray[48][84], Harray[49][84], Harray[50][84], Harray[51][84], Harray[52][84], Harray[53][84], Harray[54][84], Harray[55][84], Harray[56][84], Harray[57][84], Harray[58][84], Harray[59][84], Harray[60][84], Harray[61][84], Harray[62][84], Harray[63][84], Harray[64][84], Harray[65][84], Harray[66][84], Harray[67][84], Harray[68][84], Harray[69][84], Harray[70][84], Harray[71][84], Harray[72][84], Harray[73][84], Harray[74][84], Harray[75][84], Harray[76][84], Harray[77][84], Harray[78][84], Harray[79][84], Harray[80][84], Harray[81][84], Harray[82][84], Harray[83][84], Harray[84][84], Harray[85][84], Harray[86][84], Harray[87][84], Harray[88][84], Harray[89][84], Harray[90][84], Harray[91][84], Harray[92][84], Harray[93][84], Harray[94][84], Harray[95][84], Harray[96][84], Harray[97][84], Harray[98][84], Harray[99][84], Harray[100][84], Harray[101][84], Harray[102][84], Harray[103][84], Harray[104][84], Harray[105][84], Harray[106][84], Harray[107][84], Harray[108][84], Harray[109][84], Harray[110][84], Harray[111][84], Harray[112][84], Harray[113][84], Harray[114][84], Harray[115][84], Harray[116][84], Harray[117][84], Harray[118][84], Harray[119][84], Harray[120][84], Harray[121][84], Harray[122][84], Harray[123][84], Harray[124][84], Harray[125][84], Harray[126][84], Harray[127][84]};
assign h_col_85 = {Harray[0][85], Harray[1][85], Harray[2][85], Harray[3][85], Harray[4][85], Harray[5][85], Harray[6][85], Harray[7][85], Harray[8][85], Harray[9][85], Harray[10][85], Harray[11][85], Harray[12][85], Harray[13][85], Harray[14][85], Harray[15][85], Harray[16][85], Harray[17][85], Harray[18][85], Harray[19][85], Harray[20][85], Harray[21][85], Harray[22][85], Harray[23][85], Harray[24][85], Harray[25][85], Harray[26][85], Harray[27][85], Harray[28][85], Harray[29][85], Harray[30][85], Harray[31][85], Harray[32][85], Harray[33][85], Harray[34][85], Harray[35][85], Harray[36][85], Harray[37][85], Harray[38][85], Harray[39][85], Harray[40][85], Harray[41][85], Harray[42][85], Harray[43][85], Harray[44][85], Harray[45][85], Harray[46][85], Harray[47][85], Harray[48][85], Harray[49][85], Harray[50][85], Harray[51][85], Harray[52][85], Harray[53][85], Harray[54][85], Harray[55][85], Harray[56][85], Harray[57][85], Harray[58][85], Harray[59][85], Harray[60][85], Harray[61][85], Harray[62][85], Harray[63][85], Harray[64][85], Harray[65][85], Harray[66][85], Harray[67][85], Harray[68][85], Harray[69][85], Harray[70][85], Harray[71][85], Harray[72][85], Harray[73][85], Harray[74][85], Harray[75][85], Harray[76][85], Harray[77][85], Harray[78][85], Harray[79][85], Harray[80][85], Harray[81][85], Harray[82][85], Harray[83][85], Harray[84][85], Harray[85][85], Harray[86][85], Harray[87][85], Harray[88][85], Harray[89][85], Harray[90][85], Harray[91][85], Harray[92][85], Harray[93][85], Harray[94][85], Harray[95][85], Harray[96][85], Harray[97][85], Harray[98][85], Harray[99][85], Harray[100][85], Harray[101][85], Harray[102][85], Harray[103][85], Harray[104][85], Harray[105][85], Harray[106][85], Harray[107][85], Harray[108][85], Harray[109][85], Harray[110][85], Harray[111][85], Harray[112][85], Harray[113][85], Harray[114][85], Harray[115][85], Harray[116][85], Harray[117][85], Harray[118][85], Harray[119][85], Harray[120][85], Harray[121][85], Harray[122][85], Harray[123][85], Harray[124][85], Harray[125][85], Harray[126][85], Harray[127][85]};
assign h_col_86 = {Harray[0][86], Harray[1][86], Harray[2][86], Harray[3][86], Harray[4][86], Harray[5][86], Harray[6][86], Harray[7][86], Harray[8][86], Harray[9][86], Harray[10][86], Harray[11][86], Harray[12][86], Harray[13][86], Harray[14][86], Harray[15][86], Harray[16][86], Harray[17][86], Harray[18][86], Harray[19][86], Harray[20][86], Harray[21][86], Harray[22][86], Harray[23][86], Harray[24][86], Harray[25][86], Harray[26][86], Harray[27][86], Harray[28][86], Harray[29][86], Harray[30][86], Harray[31][86], Harray[32][86], Harray[33][86], Harray[34][86], Harray[35][86], Harray[36][86], Harray[37][86], Harray[38][86], Harray[39][86], Harray[40][86], Harray[41][86], Harray[42][86], Harray[43][86], Harray[44][86], Harray[45][86], Harray[46][86], Harray[47][86], Harray[48][86], Harray[49][86], Harray[50][86], Harray[51][86], Harray[52][86], Harray[53][86], Harray[54][86], Harray[55][86], Harray[56][86], Harray[57][86], Harray[58][86], Harray[59][86], Harray[60][86], Harray[61][86], Harray[62][86], Harray[63][86], Harray[64][86], Harray[65][86], Harray[66][86], Harray[67][86], Harray[68][86], Harray[69][86], Harray[70][86], Harray[71][86], Harray[72][86], Harray[73][86], Harray[74][86], Harray[75][86], Harray[76][86], Harray[77][86], Harray[78][86], Harray[79][86], Harray[80][86], Harray[81][86], Harray[82][86], Harray[83][86], Harray[84][86], Harray[85][86], Harray[86][86], Harray[87][86], Harray[88][86], Harray[89][86], Harray[90][86], Harray[91][86], Harray[92][86], Harray[93][86], Harray[94][86], Harray[95][86], Harray[96][86], Harray[97][86], Harray[98][86], Harray[99][86], Harray[100][86], Harray[101][86], Harray[102][86], Harray[103][86], Harray[104][86], Harray[105][86], Harray[106][86], Harray[107][86], Harray[108][86], Harray[109][86], Harray[110][86], Harray[111][86], Harray[112][86], Harray[113][86], Harray[114][86], Harray[115][86], Harray[116][86], Harray[117][86], Harray[118][86], Harray[119][86], Harray[120][86], Harray[121][86], Harray[122][86], Harray[123][86], Harray[124][86], Harray[125][86], Harray[126][86], Harray[127][86]};
assign h_col_87 = {Harray[0][87], Harray[1][87], Harray[2][87], Harray[3][87], Harray[4][87], Harray[5][87], Harray[6][87], Harray[7][87], Harray[8][87], Harray[9][87], Harray[10][87], Harray[11][87], Harray[12][87], Harray[13][87], Harray[14][87], Harray[15][87], Harray[16][87], Harray[17][87], Harray[18][87], Harray[19][87], Harray[20][87], Harray[21][87], Harray[22][87], Harray[23][87], Harray[24][87], Harray[25][87], Harray[26][87], Harray[27][87], Harray[28][87], Harray[29][87], Harray[30][87], Harray[31][87], Harray[32][87], Harray[33][87], Harray[34][87], Harray[35][87], Harray[36][87], Harray[37][87], Harray[38][87], Harray[39][87], Harray[40][87], Harray[41][87], Harray[42][87], Harray[43][87], Harray[44][87], Harray[45][87], Harray[46][87], Harray[47][87], Harray[48][87], Harray[49][87], Harray[50][87], Harray[51][87], Harray[52][87], Harray[53][87], Harray[54][87], Harray[55][87], Harray[56][87], Harray[57][87], Harray[58][87], Harray[59][87], Harray[60][87], Harray[61][87], Harray[62][87], Harray[63][87], Harray[64][87], Harray[65][87], Harray[66][87], Harray[67][87], Harray[68][87], Harray[69][87], Harray[70][87], Harray[71][87], Harray[72][87], Harray[73][87], Harray[74][87], Harray[75][87], Harray[76][87], Harray[77][87], Harray[78][87], Harray[79][87], Harray[80][87], Harray[81][87], Harray[82][87], Harray[83][87], Harray[84][87], Harray[85][87], Harray[86][87], Harray[87][87], Harray[88][87], Harray[89][87], Harray[90][87], Harray[91][87], Harray[92][87], Harray[93][87], Harray[94][87], Harray[95][87], Harray[96][87], Harray[97][87], Harray[98][87], Harray[99][87], Harray[100][87], Harray[101][87], Harray[102][87], Harray[103][87], Harray[104][87], Harray[105][87], Harray[106][87], Harray[107][87], Harray[108][87], Harray[109][87], Harray[110][87], Harray[111][87], Harray[112][87], Harray[113][87], Harray[114][87], Harray[115][87], Harray[116][87], Harray[117][87], Harray[118][87], Harray[119][87], Harray[120][87], Harray[121][87], Harray[122][87], Harray[123][87], Harray[124][87], Harray[125][87], Harray[126][87], Harray[127][87]};
assign h_col_88 = {Harray[0][88], Harray[1][88], Harray[2][88], Harray[3][88], Harray[4][88], Harray[5][88], Harray[6][88], Harray[7][88], Harray[8][88], Harray[9][88], Harray[10][88], Harray[11][88], Harray[12][88], Harray[13][88], Harray[14][88], Harray[15][88], Harray[16][88], Harray[17][88], Harray[18][88], Harray[19][88], Harray[20][88], Harray[21][88], Harray[22][88], Harray[23][88], Harray[24][88], Harray[25][88], Harray[26][88], Harray[27][88], Harray[28][88], Harray[29][88], Harray[30][88], Harray[31][88], Harray[32][88], Harray[33][88], Harray[34][88], Harray[35][88], Harray[36][88], Harray[37][88], Harray[38][88], Harray[39][88], Harray[40][88], Harray[41][88], Harray[42][88], Harray[43][88], Harray[44][88], Harray[45][88], Harray[46][88], Harray[47][88], Harray[48][88], Harray[49][88], Harray[50][88], Harray[51][88], Harray[52][88], Harray[53][88], Harray[54][88], Harray[55][88], Harray[56][88], Harray[57][88], Harray[58][88], Harray[59][88], Harray[60][88], Harray[61][88], Harray[62][88], Harray[63][88], Harray[64][88], Harray[65][88], Harray[66][88], Harray[67][88], Harray[68][88], Harray[69][88], Harray[70][88], Harray[71][88], Harray[72][88], Harray[73][88], Harray[74][88], Harray[75][88], Harray[76][88], Harray[77][88], Harray[78][88], Harray[79][88], Harray[80][88], Harray[81][88], Harray[82][88], Harray[83][88], Harray[84][88], Harray[85][88], Harray[86][88], Harray[87][88], Harray[88][88], Harray[89][88], Harray[90][88], Harray[91][88], Harray[92][88], Harray[93][88], Harray[94][88], Harray[95][88], Harray[96][88], Harray[97][88], Harray[98][88], Harray[99][88], Harray[100][88], Harray[101][88], Harray[102][88], Harray[103][88], Harray[104][88], Harray[105][88], Harray[106][88], Harray[107][88], Harray[108][88], Harray[109][88], Harray[110][88], Harray[111][88], Harray[112][88], Harray[113][88], Harray[114][88], Harray[115][88], Harray[116][88], Harray[117][88], Harray[118][88], Harray[119][88], Harray[120][88], Harray[121][88], Harray[122][88], Harray[123][88], Harray[124][88], Harray[125][88], Harray[126][88], Harray[127][88]};
assign h_col_89 = {Harray[0][89], Harray[1][89], Harray[2][89], Harray[3][89], Harray[4][89], Harray[5][89], Harray[6][89], Harray[7][89], Harray[8][89], Harray[9][89], Harray[10][89], Harray[11][89], Harray[12][89], Harray[13][89], Harray[14][89], Harray[15][89], Harray[16][89], Harray[17][89], Harray[18][89], Harray[19][89], Harray[20][89], Harray[21][89], Harray[22][89], Harray[23][89], Harray[24][89], Harray[25][89], Harray[26][89], Harray[27][89], Harray[28][89], Harray[29][89], Harray[30][89], Harray[31][89], Harray[32][89], Harray[33][89], Harray[34][89], Harray[35][89], Harray[36][89], Harray[37][89], Harray[38][89], Harray[39][89], Harray[40][89], Harray[41][89], Harray[42][89], Harray[43][89], Harray[44][89], Harray[45][89], Harray[46][89], Harray[47][89], Harray[48][89], Harray[49][89], Harray[50][89], Harray[51][89], Harray[52][89], Harray[53][89], Harray[54][89], Harray[55][89], Harray[56][89], Harray[57][89], Harray[58][89], Harray[59][89], Harray[60][89], Harray[61][89], Harray[62][89], Harray[63][89], Harray[64][89], Harray[65][89], Harray[66][89], Harray[67][89], Harray[68][89], Harray[69][89], Harray[70][89], Harray[71][89], Harray[72][89], Harray[73][89], Harray[74][89], Harray[75][89], Harray[76][89], Harray[77][89], Harray[78][89], Harray[79][89], Harray[80][89], Harray[81][89], Harray[82][89], Harray[83][89], Harray[84][89], Harray[85][89], Harray[86][89], Harray[87][89], Harray[88][89], Harray[89][89], Harray[90][89], Harray[91][89], Harray[92][89], Harray[93][89], Harray[94][89], Harray[95][89], Harray[96][89], Harray[97][89], Harray[98][89], Harray[99][89], Harray[100][89], Harray[101][89], Harray[102][89], Harray[103][89], Harray[104][89], Harray[105][89], Harray[106][89], Harray[107][89], Harray[108][89], Harray[109][89], Harray[110][89], Harray[111][89], Harray[112][89], Harray[113][89], Harray[114][89], Harray[115][89], Harray[116][89], Harray[117][89], Harray[118][89], Harray[119][89], Harray[120][89], Harray[121][89], Harray[122][89], Harray[123][89], Harray[124][89], Harray[125][89], Harray[126][89], Harray[127][89]};
assign h_col_90 = {Harray[0][90], Harray[1][90], Harray[2][90], Harray[3][90], Harray[4][90], Harray[5][90], Harray[6][90], Harray[7][90], Harray[8][90], Harray[9][90], Harray[10][90], Harray[11][90], Harray[12][90], Harray[13][90], Harray[14][90], Harray[15][90], Harray[16][90], Harray[17][90], Harray[18][90], Harray[19][90], Harray[20][90], Harray[21][90], Harray[22][90], Harray[23][90], Harray[24][90], Harray[25][90], Harray[26][90], Harray[27][90], Harray[28][90], Harray[29][90], Harray[30][90], Harray[31][90], Harray[32][90], Harray[33][90], Harray[34][90], Harray[35][90], Harray[36][90], Harray[37][90], Harray[38][90], Harray[39][90], Harray[40][90], Harray[41][90], Harray[42][90], Harray[43][90], Harray[44][90], Harray[45][90], Harray[46][90], Harray[47][90], Harray[48][90], Harray[49][90], Harray[50][90], Harray[51][90], Harray[52][90], Harray[53][90], Harray[54][90], Harray[55][90], Harray[56][90], Harray[57][90], Harray[58][90], Harray[59][90], Harray[60][90], Harray[61][90], Harray[62][90], Harray[63][90], Harray[64][90], Harray[65][90], Harray[66][90], Harray[67][90], Harray[68][90], Harray[69][90], Harray[70][90], Harray[71][90], Harray[72][90], Harray[73][90], Harray[74][90], Harray[75][90], Harray[76][90], Harray[77][90], Harray[78][90], Harray[79][90], Harray[80][90], Harray[81][90], Harray[82][90], Harray[83][90], Harray[84][90], Harray[85][90], Harray[86][90], Harray[87][90], Harray[88][90], Harray[89][90], Harray[90][90], Harray[91][90], Harray[92][90], Harray[93][90], Harray[94][90], Harray[95][90], Harray[96][90], Harray[97][90], Harray[98][90], Harray[99][90], Harray[100][90], Harray[101][90], Harray[102][90], Harray[103][90], Harray[104][90], Harray[105][90], Harray[106][90], Harray[107][90], Harray[108][90], Harray[109][90], Harray[110][90], Harray[111][90], Harray[112][90], Harray[113][90], Harray[114][90], Harray[115][90], Harray[116][90], Harray[117][90], Harray[118][90], Harray[119][90], Harray[120][90], Harray[121][90], Harray[122][90], Harray[123][90], Harray[124][90], Harray[125][90], Harray[126][90], Harray[127][90]};
assign h_col_91 = {Harray[0][91], Harray[1][91], Harray[2][91], Harray[3][91], Harray[4][91], Harray[5][91], Harray[6][91], Harray[7][91], Harray[8][91], Harray[9][91], Harray[10][91], Harray[11][91], Harray[12][91], Harray[13][91], Harray[14][91], Harray[15][91], Harray[16][91], Harray[17][91], Harray[18][91], Harray[19][91], Harray[20][91], Harray[21][91], Harray[22][91], Harray[23][91], Harray[24][91], Harray[25][91], Harray[26][91], Harray[27][91], Harray[28][91], Harray[29][91], Harray[30][91], Harray[31][91], Harray[32][91], Harray[33][91], Harray[34][91], Harray[35][91], Harray[36][91], Harray[37][91], Harray[38][91], Harray[39][91], Harray[40][91], Harray[41][91], Harray[42][91], Harray[43][91], Harray[44][91], Harray[45][91], Harray[46][91], Harray[47][91], Harray[48][91], Harray[49][91], Harray[50][91], Harray[51][91], Harray[52][91], Harray[53][91], Harray[54][91], Harray[55][91], Harray[56][91], Harray[57][91], Harray[58][91], Harray[59][91], Harray[60][91], Harray[61][91], Harray[62][91], Harray[63][91], Harray[64][91], Harray[65][91], Harray[66][91], Harray[67][91], Harray[68][91], Harray[69][91], Harray[70][91], Harray[71][91], Harray[72][91], Harray[73][91], Harray[74][91], Harray[75][91], Harray[76][91], Harray[77][91], Harray[78][91], Harray[79][91], Harray[80][91], Harray[81][91], Harray[82][91], Harray[83][91], Harray[84][91], Harray[85][91], Harray[86][91], Harray[87][91], Harray[88][91], Harray[89][91], Harray[90][91], Harray[91][91], Harray[92][91], Harray[93][91], Harray[94][91], Harray[95][91], Harray[96][91], Harray[97][91], Harray[98][91], Harray[99][91], Harray[100][91], Harray[101][91], Harray[102][91], Harray[103][91], Harray[104][91], Harray[105][91], Harray[106][91], Harray[107][91], Harray[108][91], Harray[109][91], Harray[110][91], Harray[111][91], Harray[112][91], Harray[113][91], Harray[114][91], Harray[115][91], Harray[116][91], Harray[117][91], Harray[118][91], Harray[119][91], Harray[120][91], Harray[121][91], Harray[122][91], Harray[123][91], Harray[124][91], Harray[125][91], Harray[126][91], Harray[127][91]};
assign h_col_92 = {Harray[0][92], Harray[1][92], Harray[2][92], Harray[3][92], Harray[4][92], Harray[5][92], Harray[6][92], Harray[7][92], Harray[8][92], Harray[9][92], Harray[10][92], Harray[11][92], Harray[12][92], Harray[13][92], Harray[14][92], Harray[15][92], Harray[16][92], Harray[17][92], Harray[18][92], Harray[19][92], Harray[20][92], Harray[21][92], Harray[22][92], Harray[23][92], Harray[24][92], Harray[25][92], Harray[26][92], Harray[27][92], Harray[28][92], Harray[29][92], Harray[30][92], Harray[31][92], Harray[32][92], Harray[33][92], Harray[34][92], Harray[35][92], Harray[36][92], Harray[37][92], Harray[38][92], Harray[39][92], Harray[40][92], Harray[41][92], Harray[42][92], Harray[43][92], Harray[44][92], Harray[45][92], Harray[46][92], Harray[47][92], Harray[48][92], Harray[49][92], Harray[50][92], Harray[51][92], Harray[52][92], Harray[53][92], Harray[54][92], Harray[55][92], Harray[56][92], Harray[57][92], Harray[58][92], Harray[59][92], Harray[60][92], Harray[61][92], Harray[62][92], Harray[63][92], Harray[64][92], Harray[65][92], Harray[66][92], Harray[67][92], Harray[68][92], Harray[69][92], Harray[70][92], Harray[71][92], Harray[72][92], Harray[73][92], Harray[74][92], Harray[75][92], Harray[76][92], Harray[77][92], Harray[78][92], Harray[79][92], Harray[80][92], Harray[81][92], Harray[82][92], Harray[83][92], Harray[84][92], Harray[85][92], Harray[86][92], Harray[87][92], Harray[88][92], Harray[89][92], Harray[90][92], Harray[91][92], Harray[92][92], Harray[93][92], Harray[94][92], Harray[95][92], Harray[96][92], Harray[97][92], Harray[98][92], Harray[99][92], Harray[100][92], Harray[101][92], Harray[102][92], Harray[103][92], Harray[104][92], Harray[105][92], Harray[106][92], Harray[107][92], Harray[108][92], Harray[109][92], Harray[110][92], Harray[111][92], Harray[112][92], Harray[113][92], Harray[114][92], Harray[115][92], Harray[116][92], Harray[117][92], Harray[118][92], Harray[119][92], Harray[120][92], Harray[121][92], Harray[122][92], Harray[123][92], Harray[124][92], Harray[125][92], Harray[126][92], Harray[127][92]};
assign h_col_93 = {Harray[0][93], Harray[1][93], Harray[2][93], Harray[3][93], Harray[4][93], Harray[5][93], Harray[6][93], Harray[7][93], Harray[8][93], Harray[9][93], Harray[10][93], Harray[11][93], Harray[12][93], Harray[13][93], Harray[14][93], Harray[15][93], Harray[16][93], Harray[17][93], Harray[18][93], Harray[19][93], Harray[20][93], Harray[21][93], Harray[22][93], Harray[23][93], Harray[24][93], Harray[25][93], Harray[26][93], Harray[27][93], Harray[28][93], Harray[29][93], Harray[30][93], Harray[31][93], Harray[32][93], Harray[33][93], Harray[34][93], Harray[35][93], Harray[36][93], Harray[37][93], Harray[38][93], Harray[39][93], Harray[40][93], Harray[41][93], Harray[42][93], Harray[43][93], Harray[44][93], Harray[45][93], Harray[46][93], Harray[47][93], Harray[48][93], Harray[49][93], Harray[50][93], Harray[51][93], Harray[52][93], Harray[53][93], Harray[54][93], Harray[55][93], Harray[56][93], Harray[57][93], Harray[58][93], Harray[59][93], Harray[60][93], Harray[61][93], Harray[62][93], Harray[63][93], Harray[64][93], Harray[65][93], Harray[66][93], Harray[67][93], Harray[68][93], Harray[69][93], Harray[70][93], Harray[71][93], Harray[72][93], Harray[73][93], Harray[74][93], Harray[75][93], Harray[76][93], Harray[77][93], Harray[78][93], Harray[79][93], Harray[80][93], Harray[81][93], Harray[82][93], Harray[83][93], Harray[84][93], Harray[85][93], Harray[86][93], Harray[87][93], Harray[88][93], Harray[89][93], Harray[90][93], Harray[91][93], Harray[92][93], Harray[93][93], Harray[94][93], Harray[95][93], Harray[96][93], Harray[97][93], Harray[98][93], Harray[99][93], Harray[100][93], Harray[101][93], Harray[102][93], Harray[103][93], Harray[104][93], Harray[105][93], Harray[106][93], Harray[107][93], Harray[108][93], Harray[109][93], Harray[110][93], Harray[111][93], Harray[112][93], Harray[113][93], Harray[114][93], Harray[115][93], Harray[116][93], Harray[117][93], Harray[118][93], Harray[119][93], Harray[120][93], Harray[121][93], Harray[122][93], Harray[123][93], Harray[124][93], Harray[125][93], Harray[126][93], Harray[127][93]};
assign h_col_94 = {Harray[0][94], Harray[1][94], Harray[2][94], Harray[3][94], Harray[4][94], Harray[5][94], Harray[6][94], Harray[7][94], Harray[8][94], Harray[9][94], Harray[10][94], Harray[11][94], Harray[12][94], Harray[13][94], Harray[14][94], Harray[15][94], Harray[16][94], Harray[17][94], Harray[18][94], Harray[19][94], Harray[20][94], Harray[21][94], Harray[22][94], Harray[23][94], Harray[24][94], Harray[25][94], Harray[26][94], Harray[27][94], Harray[28][94], Harray[29][94], Harray[30][94], Harray[31][94], Harray[32][94], Harray[33][94], Harray[34][94], Harray[35][94], Harray[36][94], Harray[37][94], Harray[38][94], Harray[39][94], Harray[40][94], Harray[41][94], Harray[42][94], Harray[43][94], Harray[44][94], Harray[45][94], Harray[46][94], Harray[47][94], Harray[48][94], Harray[49][94], Harray[50][94], Harray[51][94], Harray[52][94], Harray[53][94], Harray[54][94], Harray[55][94], Harray[56][94], Harray[57][94], Harray[58][94], Harray[59][94], Harray[60][94], Harray[61][94], Harray[62][94], Harray[63][94], Harray[64][94], Harray[65][94], Harray[66][94], Harray[67][94], Harray[68][94], Harray[69][94], Harray[70][94], Harray[71][94], Harray[72][94], Harray[73][94], Harray[74][94], Harray[75][94], Harray[76][94], Harray[77][94], Harray[78][94], Harray[79][94], Harray[80][94], Harray[81][94], Harray[82][94], Harray[83][94], Harray[84][94], Harray[85][94], Harray[86][94], Harray[87][94], Harray[88][94], Harray[89][94], Harray[90][94], Harray[91][94], Harray[92][94], Harray[93][94], Harray[94][94], Harray[95][94], Harray[96][94], Harray[97][94], Harray[98][94], Harray[99][94], Harray[100][94], Harray[101][94], Harray[102][94], Harray[103][94], Harray[104][94], Harray[105][94], Harray[106][94], Harray[107][94], Harray[108][94], Harray[109][94], Harray[110][94], Harray[111][94], Harray[112][94], Harray[113][94], Harray[114][94], Harray[115][94], Harray[116][94], Harray[117][94], Harray[118][94], Harray[119][94], Harray[120][94], Harray[121][94], Harray[122][94], Harray[123][94], Harray[124][94], Harray[125][94], Harray[126][94], Harray[127][94]};
assign h_col_95 = {Harray[0][95], Harray[1][95], Harray[2][95], Harray[3][95], Harray[4][95], Harray[5][95], Harray[6][95], Harray[7][95], Harray[8][95], Harray[9][95], Harray[10][95], Harray[11][95], Harray[12][95], Harray[13][95], Harray[14][95], Harray[15][95], Harray[16][95], Harray[17][95], Harray[18][95], Harray[19][95], Harray[20][95], Harray[21][95], Harray[22][95], Harray[23][95], Harray[24][95], Harray[25][95], Harray[26][95], Harray[27][95], Harray[28][95], Harray[29][95], Harray[30][95], Harray[31][95], Harray[32][95], Harray[33][95], Harray[34][95], Harray[35][95], Harray[36][95], Harray[37][95], Harray[38][95], Harray[39][95], Harray[40][95], Harray[41][95], Harray[42][95], Harray[43][95], Harray[44][95], Harray[45][95], Harray[46][95], Harray[47][95], Harray[48][95], Harray[49][95], Harray[50][95], Harray[51][95], Harray[52][95], Harray[53][95], Harray[54][95], Harray[55][95], Harray[56][95], Harray[57][95], Harray[58][95], Harray[59][95], Harray[60][95], Harray[61][95], Harray[62][95], Harray[63][95], Harray[64][95], Harray[65][95], Harray[66][95], Harray[67][95], Harray[68][95], Harray[69][95], Harray[70][95], Harray[71][95], Harray[72][95], Harray[73][95], Harray[74][95], Harray[75][95], Harray[76][95], Harray[77][95], Harray[78][95], Harray[79][95], Harray[80][95], Harray[81][95], Harray[82][95], Harray[83][95], Harray[84][95], Harray[85][95], Harray[86][95], Harray[87][95], Harray[88][95], Harray[89][95], Harray[90][95], Harray[91][95], Harray[92][95], Harray[93][95], Harray[94][95], Harray[95][95], Harray[96][95], Harray[97][95], Harray[98][95], Harray[99][95], Harray[100][95], Harray[101][95], Harray[102][95], Harray[103][95], Harray[104][95], Harray[105][95], Harray[106][95], Harray[107][95], Harray[108][95], Harray[109][95], Harray[110][95], Harray[111][95], Harray[112][95], Harray[113][95], Harray[114][95], Harray[115][95], Harray[116][95], Harray[117][95], Harray[118][95], Harray[119][95], Harray[120][95], Harray[121][95], Harray[122][95], Harray[123][95], Harray[124][95], Harray[125][95], Harray[126][95], Harray[127][95]};
assign h_col_96 = {Harray[0][96], Harray[1][96], Harray[2][96], Harray[3][96], Harray[4][96], Harray[5][96], Harray[6][96], Harray[7][96], Harray[8][96], Harray[9][96], Harray[10][96], Harray[11][96], Harray[12][96], Harray[13][96], Harray[14][96], Harray[15][96], Harray[16][96], Harray[17][96], Harray[18][96], Harray[19][96], Harray[20][96], Harray[21][96], Harray[22][96], Harray[23][96], Harray[24][96], Harray[25][96], Harray[26][96], Harray[27][96], Harray[28][96], Harray[29][96], Harray[30][96], Harray[31][96], Harray[32][96], Harray[33][96], Harray[34][96], Harray[35][96], Harray[36][96], Harray[37][96], Harray[38][96], Harray[39][96], Harray[40][96], Harray[41][96], Harray[42][96], Harray[43][96], Harray[44][96], Harray[45][96], Harray[46][96], Harray[47][96], Harray[48][96], Harray[49][96], Harray[50][96], Harray[51][96], Harray[52][96], Harray[53][96], Harray[54][96], Harray[55][96], Harray[56][96], Harray[57][96], Harray[58][96], Harray[59][96], Harray[60][96], Harray[61][96], Harray[62][96], Harray[63][96], Harray[64][96], Harray[65][96], Harray[66][96], Harray[67][96], Harray[68][96], Harray[69][96], Harray[70][96], Harray[71][96], Harray[72][96], Harray[73][96], Harray[74][96], Harray[75][96], Harray[76][96], Harray[77][96], Harray[78][96], Harray[79][96], Harray[80][96], Harray[81][96], Harray[82][96], Harray[83][96], Harray[84][96], Harray[85][96], Harray[86][96], Harray[87][96], Harray[88][96], Harray[89][96], Harray[90][96], Harray[91][96], Harray[92][96], Harray[93][96], Harray[94][96], Harray[95][96], Harray[96][96], Harray[97][96], Harray[98][96], Harray[99][96], Harray[100][96], Harray[101][96], Harray[102][96], Harray[103][96], Harray[104][96], Harray[105][96], Harray[106][96], Harray[107][96], Harray[108][96], Harray[109][96], Harray[110][96], Harray[111][96], Harray[112][96], Harray[113][96], Harray[114][96], Harray[115][96], Harray[116][96], Harray[117][96], Harray[118][96], Harray[119][96], Harray[120][96], Harray[121][96], Harray[122][96], Harray[123][96], Harray[124][96], Harray[125][96], Harray[126][96], Harray[127][96]};
assign h_col_97 = {Harray[0][97], Harray[1][97], Harray[2][97], Harray[3][97], Harray[4][97], Harray[5][97], Harray[6][97], Harray[7][97], Harray[8][97], Harray[9][97], Harray[10][97], Harray[11][97], Harray[12][97], Harray[13][97], Harray[14][97], Harray[15][97], Harray[16][97], Harray[17][97], Harray[18][97], Harray[19][97], Harray[20][97], Harray[21][97], Harray[22][97], Harray[23][97], Harray[24][97], Harray[25][97], Harray[26][97], Harray[27][97], Harray[28][97], Harray[29][97], Harray[30][97], Harray[31][97], Harray[32][97], Harray[33][97], Harray[34][97], Harray[35][97], Harray[36][97], Harray[37][97], Harray[38][97], Harray[39][97], Harray[40][97], Harray[41][97], Harray[42][97], Harray[43][97], Harray[44][97], Harray[45][97], Harray[46][97], Harray[47][97], Harray[48][97], Harray[49][97], Harray[50][97], Harray[51][97], Harray[52][97], Harray[53][97], Harray[54][97], Harray[55][97], Harray[56][97], Harray[57][97], Harray[58][97], Harray[59][97], Harray[60][97], Harray[61][97], Harray[62][97], Harray[63][97], Harray[64][97], Harray[65][97], Harray[66][97], Harray[67][97], Harray[68][97], Harray[69][97], Harray[70][97], Harray[71][97], Harray[72][97], Harray[73][97], Harray[74][97], Harray[75][97], Harray[76][97], Harray[77][97], Harray[78][97], Harray[79][97], Harray[80][97], Harray[81][97], Harray[82][97], Harray[83][97], Harray[84][97], Harray[85][97], Harray[86][97], Harray[87][97], Harray[88][97], Harray[89][97], Harray[90][97], Harray[91][97], Harray[92][97], Harray[93][97], Harray[94][97], Harray[95][97], Harray[96][97], Harray[97][97], Harray[98][97], Harray[99][97], Harray[100][97], Harray[101][97], Harray[102][97], Harray[103][97], Harray[104][97], Harray[105][97], Harray[106][97], Harray[107][97], Harray[108][97], Harray[109][97], Harray[110][97], Harray[111][97], Harray[112][97], Harray[113][97], Harray[114][97], Harray[115][97], Harray[116][97], Harray[117][97], Harray[118][97], Harray[119][97], Harray[120][97], Harray[121][97], Harray[122][97], Harray[123][97], Harray[124][97], Harray[125][97], Harray[126][97], Harray[127][97]};
assign h_col_98 = {Harray[0][98], Harray[1][98], Harray[2][98], Harray[3][98], Harray[4][98], Harray[5][98], Harray[6][98], Harray[7][98], Harray[8][98], Harray[9][98], Harray[10][98], Harray[11][98], Harray[12][98], Harray[13][98], Harray[14][98], Harray[15][98], Harray[16][98], Harray[17][98], Harray[18][98], Harray[19][98], Harray[20][98], Harray[21][98], Harray[22][98], Harray[23][98], Harray[24][98], Harray[25][98], Harray[26][98], Harray[27][98], Harray[28][98], Harray[29][98], Harray[30][98], Harray[31][98], Harray[32][98], Harray[33][98], Harray[34][98], Harray[35][98], Harray[36][98], Harray[37][98], Harray[38][98], Harray[39][98], Harray[40][98], Harray[41][98], Harray[42][98], Harray[43][98], Harray[44][98], Harray[45][98], Harray[46][98], Harray[47][98], Harray[48][98], Harray[49][98], Harray[50][98], Harray[51][98], Harray[52][98], Harray[53][98], Harray[54][98], Harray[55][98], Harray[56][98], Harray[57][98], Harray[58][98], Harray[59][98], Harray[60][98], Harray[61][98], Harray[62][98], Harray[63][98], Harray[64][98], Harray[65][98], Harray[66][98], Harray[67][98], Harray[68][98], Harray[69][98], Harray[70][98], Harray[71][98], Harray[72][98], Harray[73][98], Harray[74][98], Harray[75][98], Harray[76][98], Harray[77][98], Harray[78][98], Harray[79][98], Harray[80][98], Harray[81][98], Harray[82][98], Harray[83][98], Harray[84][98], Harray[85][98], Harray[86][98], Harray[87][98], Harray[88][98], Harray[89][98], Harray[90][98], Harray[91][98], Harray[92][98], Harray[93][98], Harray[94][98], Harray[95][98], Harray[96][98], Harray[97][98], Harray[98][98], Harray[99][98], Harray[100][98], Harray[101][98], Harray[102][98], Harray[103][98], Harray[104][98], Harray[105][98], Harray[106][98], Harray[107][98], Harray[108][98], Harray[109][98], Harray[110][98], Harray[111][98], Harray[112][98], Harray[113][98], Harray[114][98], Harray[115][98], Harray[116][98], Harray[117][98], Harray[118][98], Harray[119][98], Harray[120][98], Harray[121][98], Harray[122][98], Harray[123][98], Harray[124][98], Harray[125][98], Harray[126][98], Harray[127][98]};
assign h_col_99 = {Harray[0][99], Harray[1][99], Harray[2][99], Harray[3][99], Harray[4][99], Harray[5][99], Harray[6][99], Harray[7][99], Harray[8][99], Harray[9][99], Harray[10][99], Harray[11][99], Harray[12][99], Harray[13][99], Harray[14][99], Harray[15][99], Harray[16][99], Harray[17][99], Harray[18][99], Harray[19][99], Harray[20][99], Harray[21][99], Harray[22][99], Harray[23][99], Harray[24][99], Harray[25][99], Harray[26][99], Harray[27][99], Harray[28][99], Harray[29][99], Harray[30][99], Harray[31][99], Harray[32][99], Harray[33][99], Harray[34][99], Harray[35][99], Harray[36][99], Harray[37][99], Harray[38][99], Harray[39][99], Harray[40][99], Harray[41][99], Harray[42][99], Harray[43][99], Harray[44][99], Harray[45][99], Harray[46][99], Harray[47][99], Harray[48][99], Harray[49][99], Harray[50][99], Harray[51][99], Harray[52][99], Harray[53][99], Harray[54][99], Harray[55][99], Harray[56][99], Harray[57][99], Harray[58][99], Harray[59][99], Harray[60][99], Harray[61][99], Harray[62][99], Harray[63][99], Harray[64][99], Harray[65][99], Harray[66][99], Harray[67][99], Harray[68][99], Harray[69][99], Harray[70][99], Harray[71][99], Harray[72][99], Harray[73][99], Harray[74][99], Harray[75][99], Harray[76][99], Harray[77][99], Harray[78][99], Harray[79][99], Harray[80][99], Harray[81][99], Harray[82][99], Harray[83][99], Harray[84][99], Harray[85][99], Harray[86][99], Harray[87][99], Harray[88][99], Harray[89][99], Harray[90][99], Harray[91][99], Harray[92][99], Harray[93][99], Harray[94][99], Harray[95][99], Harray[96][99], Harray[97][99], Harray[98][99], Harray[99][99], Harray[100][99], Harray[101][99], Harray[102][99], Harray[103][99], Harray[104][99], Harray[105][99], Harray[106][99], Harray[107][99], Harray[108][99], Harray[109][99], Harray[110][99], Harray[111][99], Harray[112][99], Harray[113][99], Harray[114][99], Harray[115][99], Harray[116][99], Harray[117][99], Harray[118][99], Harray[119][99], Harray[120][99], Harray[121][99], Harray[122][99], Harray[123][99], Harray[124][99], Harray[125][99], Harray[126][99], Harray[127][99]};
assign h_col_100 = {Harray[0][100], Harray[1][100], Harray[2][100], Harray[3][100], Harray[4][100], Harray[5][100], Harray[6][100], Harray[7][100], Harray[8][100], Harray[9][100], Harray[10][100], Harray[11][100], Harray[12][100], Harray[13][100], Harray[14][100], Harray[15][100], Harray[16][100], Harray[17][100], Harray[18][100], Harray[19][100], Harray[20][100], Harray[21][100], Harray[22][100], Harray[23][100], Harray[24][100], Harray[25][100], Harray[26][100], Harray[27][100], Harray[28][100], Harray[29][100], Harray[30][100], Harray[31][100], Harray[32][100], Harray[33][100], Harray[34][100], Harray[35][100], Harray[36][100], Harray[37][100], Harray[38][100], Harray[39][100], Harray[40][100], Harray[41][100], Harray[42][100], Harray[43][100], Harray[44][100], Harray[45][100], Harray[46][100], Harray[47][100], Harray[48][100], Harray[49][100], Harray[50][100], Harray[51][100], Harray[52][100], Harray[53][100], Harray[54][100], Harray[55][100], Harray[56][100], Harray[57][100], Harray[58][100], Harray[59][100], Harray[60][100], Harray[61][100], Harray[62][100], Harray[63][100], Harray[64][100], Harray[65][100], Harray[66][100], Harray[67][100], Harray[68][100], Harray[69][100], Harray[70][100], Harray[71][100], Harray[72][100], Harray[73][100], Harray[74][100], Harray[75][100], Harray[76][100], Harray[77][100], Harray[78][100], Harray[79][100], Harray[80][100], Harray[81][100], Harray[82][100], Harray[83][100], Harray[84][100], Harray[85][100], Harray[86][100], Harray[87][100], Harray[88][100], Harray[89][100], Harray[90][100], Harray[91][100], Harray[92][100], Harray[93][100], Harray[94][100], Harray[95][100], Harray[96][100], Harray[97][100], Harray[98][100], Harray[99][100], Harray[100][100], Harray[101][100], Harray[102][100], Harray[103][100], Harray[104][100], Harray[105][100], Harray[106][100], Harray[107][100], Harray[108][100], Harray[109][100], Harray[110][100], Harray[111][100], Harray[112][100], Harray[113][100], Harray[114][100], Harray[115][100], Harray[116][100], Harray[117][100], Harray[118][100], Harray[119][100], Harray[120][100], Harray[121][100], Harray[122][100], Harray[123][100], Harray[124][100], Harray[125][100], Harray[126][100], Harray[127][100]};
assign h_col_101 = {Harray[0][101], Harray[1][101], Harray[2][101], Harray[3][101], Harray[4][101], Harray[5][101], Harray[6][101], Harray[7][101], Harray[8][101], Harray[9][101], Harray[10][101], Harray[11][101], Harray[12][101], Harray[13][101], Harray[14][101], Harray[15][101], Harray[16][101], Harray[17][101], Harray[18][101], Harray[19][101], Harray[20][101], Harray[21][101], Harray[22][101], Harray[23][101], Harray[24][101], Harray[25][101], Harray[26][101], Harray[27][101], Harray[28][101], Harray[29][101], Harray[30][101], Harray[31][101], Harray[32][101], Harray[33][101], Harray[34][101], Harray[35][101], Harray[36][101], Harray[37][101], Harray[38][101], Harray[39][101], Harray[40][101], Harray[41][101], Harray[42][101], Harray[43][101], Harray[44][101], Harray[45][101], Harray[46][101], Harray[47][101], Harray[48][101], Harray[49][101], Harray[50][101], Harray[51][101], Harray[52][101], Harray[53][101], Harray[54][101], Harray[55][101], Harray[56][101], Harray[57][101], Harray[58][101], Harray[59][101], Harray[60][101], Harray[61][101], Harray[62][101], Harray[63][101], Harray[64][101], Harray[65][101], Harray[66][101], Harray[67][101], Harray[68][101], Harray[69][101], Harray[70][101], Harray[71][101], Harray[72][101], Harray[73][101], Harray[74][101], Harray[75][101], Harray[76][101], Harray[77][101], Harray[78][101], Harray[79][101], Harray[80][101], Harray[81][101], Harray[82][101], Harray[83][101], Harray[84][101], Harray[85][101], Harray[86][101], Harray[87][101], Harray[88][101], Harray[89][101], Harray[90][101], Harray[91][101], Harray[92][101], Harray[93][101], Harray[94][101], Harray[95][101], Harray[96][101], Harray[97][101], Harray[98][101], Harray[99][101], Harray[100][101], Harray[101][101], Harray[102][101], Harray[103][101], Harray[104][101], Harray[105][101], Harray[106][101], Harray[107][101], Harray[108][101], Harray[109][101], Harray[110][101], Harray[111][101], Harray[112][101], Harray[113][101], Harray[114][101], Harray[115][101], Harray[116][101], Harray[117][101], Harray[118][101], Harray[119][101], Harray[120][101], Harray[121][101], Harray[122][101], Harray[123][101], Harray[124][101], Harray[125][101], Harray[126][101], Harray[127][101]};
assign h_col_102 = {Harray[0][102], Harray[1][102], Harray[2][102], Harray[3][102], Harray[4][102], Harray[5][102], Harray[6][102], Harray[7][102], Harray[8][102], Harray[9][102], Harray[10][102], Harray[11][102], Harray[12][102], Harray[13][102], Harray[14][102], Harray[15][102], Harray[16][102], Harray[17][102], Harray[18][102], Harray[19][102], Harray[20][102], Harray[21][102], Harray[22][102], Harray[23][102], Harray[24][102], Harray[25][102], Harray[26][102], Harray[27][102], Harray[28][102], Harray[29][102], Harray[30][102], Harray[31][102], Harray[32][102], Harray[33][102], Harray[34][102], Harray[35][102], Harray[36][102], Harray[37][102], Harray[38][102], Harray[39][102], Harray[40][102], Harray[41][102], Harray[42][102], Harray[43][102], Harray[44][102], Harray[45][102], Harray[46][102], Harray[47][102], Harray[48][102], Harray[49][102], Harray[50][102], Harray[51][102], Harray[52][102], Harray[53][102], Harray[54][102], Harray[55][102], Harray[56][102], Harray[57][102], Harray[58][102], Harray[59][102], Harray[60][102], Harray[61][102], Harray[62][102], Harray[63][102], Harray[64][102], Harray[65][102], Harray[66][102], Harray[67][102], Harray[68][102], Harray[69][102], Harray[70][102], Harray[71][102], Harray[72][102], Harray[73][102], Harray[74][102], Harray[75][102], Harray[76][102], Harray[77][102], Harray[78][102], Harray[79][102], Harray[80][102], Harray[81][102], Harray[82][102], Harray[83][102], Harray[84][102], Harray[85][102], Harray[86][102], Harray[87][102], Harray[88][102], Harray[89][102], Harray[90][102], Harray[91][102], Harray[92][102], Harray[93][102], Harray[94][102], Harray[95][102], Harray[96][102], Harray[97][102], Harray[98][102], Harray[99][102], Harray[100][102], Harray[101][102], Harray[102][102], Harray[103][102], Harray[104][102], Harray[105][102], Harray[106][102], Harray[107][102], Harray[108][102], Harray[109][102], Harray[110][102], Harray[111][102], Harray[112][102], Harray[113][102], Harray[114][102], Harray[115][102], Harray[116][102], Harray[117][102], Harray[118][102], Harray[119][102], Harray[120][102], Harray[121][102], Harray[122][102], Harray[123][102], Harray[124][102], Harray[125][102], Harray[126][102], Harray[127][102]};
assign h_col_103 = {Harray[0][103], Harray[1][103], Harray[2][103], Harray[3][103], Harray[4][103], Harray[5][103], Harray[6][103], Harray[7][103], Harray[8][103], Harray[9][103], Harray[10][103], Harray[11][103], Harray[12][103], Harray[13][103], Harray[14][103], Harray[15][103], Harray[16][103], Harray[17][103], Harray[18][103], Harray[19][103], Harray[20][103], Harray[21][103], Harray[22][103], Harray[23][103], Harray[24][103], Harray[25][103], Harray[26][103], Harray[27][103], Harray[28][103], Harray[29][103], Harray[30][103], Harray[31][103], Harray[32][103], Harray[33][103], Harray[34][103], Harray[35][103], Harray[36][103], Harray[37][103], Harray[38][103], Harray[39][103], Harray[40][103], Harray[41][103], Harray[42][103], Harray[43][103], Harray[44][103], Harray[45][103], Harray[46][103], Harray[47][103], Harray[48][103], Harray[49][103], Harray[50][103], Harray[51][103], Harray[52][103], Harray[53][103], Harray[54][103], Harray[55][103], Harray[56][103], Harray[57][103], Harray[58][103], Harray[59][103], Harray[60][103], Harray[61][103], Harray[62][103], Harray[63][103], Harray[64][103], Harray[65][103], Harray[66][103], Harray[67][103], Harray[68][103], Harray[69][103], Harray[70][103], Harray[71][103], Harray[72][103], Harray[73][103], Harray[74][103], Harray[75][103], Harray[76][103], Harray[77][103], Harray[78][103], Harray[79][103], Harray[80][103], Harray[81][103], Harray[82][103], Harray[83][103], Harray[84][103], Harray[85][103], Harray[86][103], Harray[87][103], Harray[88][103], Harray[89][103], Harray[90][103], Harray[91][103], Harray[92][103], Harray[93][103], Harray[94][103], Harray[95][103], Harray[96][103], Harray[97][103], Harray[98][103], Harray[99][103], Harray[100][103], Harray[101][103], Harray[102][103], Harray[103][103], Harray[104][103], Harray[105][103], Harray[106][103], Harray[107][103], Harray[108][103], Harray[109][103], Harray[110][103], Harray[111][103], Harray[112][103], Harray[113][103], Harray[114][103], Harray[115][103], Harray[116][103], Harray[117][103], Harray[118][103], Harray[119][103], Harray[120][103], Harray[121][103], Harray[122][103], Harray[123][103], Harray[124][103], Harray[125][103], Harray[126][103], Harray[127][103]};
assign h_col_104 = {Harray[0][104], Harray[1][104], Harray[2][104], Harray[3][104], Harray[4][104], Harray[5][104], Harray[6][104], Harray[7][104], Harray[8][104], Harray[9][104], Harray[10][104], Harray[11][104], Harray[12][104], Harray[13][104], Harray[14][104], Harray[15][104], Harray[16][104], Harray[17][104], Harray[18][104], Harray[19][104], Harray[20][104], Harray[21][104], Harray[22][104], Harray[23][104], Harray[24][104], Harray[25][104], Harray[26][104], Harray[27][104], Harray[28][104], Harray[29][104], Harray[30][104], Harray[31][104], Harray[32][104], Harray[33][104], Harray[34][104], Harray[35][104], Harray[36][104], Harray[37][104], Harray[38][104], Harray[39][104], Harray[40][104], Harray[41][104], Harray[42][104], Harray[43][104], Harray[44][104], Harray[45][104], Harray[46][104], Harray[47][104], Harray[48][104], Harray[49][104], Harray[50][104], Harray[51][104], Harray[52][104], Harray[53][104], Harray[54][104], Harray[55][104], Harray[56][104], Harray[57][104], Harray[58][104], Harray[59][104], Harray[60][104], Harray[61][104], Harray[62][104], Harray[63][104], Harray[64][104], Harray[65][104], Harray[66][104], Harray[67][104], Harray[68][104], Harray[69][104], Harray[70][104], Harray[71][104], Harray[72][104], Harray[73][104], Harray[74][104], Harray[75][104], Harray[76][104], Harray[77][104], Harray[78][104], Harray[79][104], Harray[80][104], Harray[81][104], Harray[82][104], Harray[83][104], Harray[84][104], Harray[85][104], Harray[86][104], Harray[87][104], Harray[88][104], Harray[89][104], Harray[90][104], Harray[91][104], Harray[92][104], Harray[93][104], Harray[94][104], Harray[95][104], Harray[96][104], Harray[97][104], Harray[98][104], Harray[99][104], Harray[100][104], Harray[101][104], Harray[102][104], Harray[103][104], Harray[104][104], Harray[105][104], Harray[106][104], Harray[107][104], Harray[108][104], Harray[109][104], Harray[110][104], Harray[111][104], Harray[112][104], Harray[113][104], Harray[114][104], Harray[115][104], Harray[116][104], Harray[117][104], Harray[118][104], Harray[119][104], Harray[120][104], Harray[121][104], Harray[122][104], Harray[123][104], Harray[124][104], Harray[125][104], Harray[126][104], Harray[127][104]};
assign h_col_105 = {Harray[0][105], Harray[1][105], Harray[2][105], Harray[3][105], Harray[4][105], Harray[5][105], Harray[6][105], Harray[7][105], Harray[8][105], Harray[9][105], Harray[10][105], Harray[11][105], Harray[12][105], Harray[13][105], Harray[14][105], Harray[15][105], Harray[16][105], Harray[17][105], Harray[18][105], Harray[19][105], Harray[20][105], Harray[21][105], Harray[22][105], Harray[23][105], Harray[24][105], Harray[25][105], Harray[26][105], Harray[27][105], Harray[28][105], Harray[29][105], Harray[30][105], Harray[31][105], Harray[32][105], Harray[33][105], Harray[34][105], Harray[35][105], Harray[36][105], Harray[37][105], Harray[38][105], Harray[39][105], Harray[40][105], Harray[41][105], Harray[42][105], Harray[43][105], Harray[44][105], Harray[45][105], Harray[46][105], Harray[47][105], Harray[48][105], Harray[49][105], Harray[50][105], Harray[51][105], Harray[52][105], Harray[53][105], Harray[54][105], Harray[55][105], Harray[56][105], Harray[57][105], Harray[58][105], Harray[59][105], Harray[60][105], Harray[61][105], Harray[62][105], Harray[63][105], Harray[64][105], Harray[65][105], Harray[66][105], Harray[67][105], Harray[68][105], Harray[69][105], Harray[70][105], Harray[71][105], Harray[72][105], Harray[73][105], Harray[74][105], Harray[75][105], Harray[76][105], Harray[77][105], Harray[78][105], Harray[79][105], Harray[80][105], Harray[81][105], Harray[82][105], Harray[83][105], Harray[84][105], Harray[85][105], Harray[86][105], Harray[87][105], Harray[88][105], Harray[89][105], Harray[90][105], Harray[91][105], Harray[92][105], Harray[93][105], Harray[94][105], Harray[95][105], Harray[96][105], Harray[97][105], Harray[98][105], Harray[99][105], Harray[100][105], Harray[101][105], Harray[102][105], Harray[103][105], Harray[104][105], Harray[105][105], Harray[106][105], Harray[107][105], Harray[108][105], Harray[109][105], Harray[110][105], Harray[111][105], Harray[112][105], Harray[113][105], Harray[114][105], Harray[115][105], Harray[116][105], Harray[117][105], Harray[118][105], Harray[119][105], Harray[120][105], Harray[121][105], Harray[122][105], Harray[123][105], Harray[124][105], Harray[125][105], Harray[126][105], Harray[127][105]};
assign h_col_106 = {Harray[0][106], Harray[1][106], Harray[2][106], Harray[3][106], Harray[4][106], Harray[5][106], Harray[6][106], Harray[7][106], Harray[8][106], Harray[9][106], Harray[10][106], Harray[11][106], Harray[12][106], Harray[13][106], Harray[14][106], Harray[15][106], Harray[16][106], Harray[17][106], Harray[18][106], Harray[19][106], Harray[20][106], Harray[21][106], Harray[22][106], Harray[23][106], Harray[24][106], Harray[25][106], Harray[26][106], Harray[27][106], Harray[28][106], Harray[29][106], Harray[30][106], Harray[31][106], Harray[32][106], Harray[33][106], Harray[34][106], Harray[35][106], Harray[36][106], Harray[37][106], Harray[38][106], Harray[39][106], Harray[40][106], Harray[41][106], Harray[42][106], Harray[43][106], Harray[44][106], Harray[45][106], Harray[46][106], Harray[47][106], Harray[48][106], Harray[49][106], Harray[50][106], Harray[51][106], Harray[52][106], Harray[53][106], Harray[54][106], Harray[55][106], Harray[56][106], Harray[57][106], Harray[58][106], Harray[59][106], Harray[60][106], Harray[61][106], Harray[62][106], Harray[63][106], Harray[64][106], Harray[65][106], Harray[66][106], Harray[67][106], Harray[68][106], Harray[69][106], Harray[70][106], Harray[71][106], Harray[72][106], Harray[73][106], Harray[74][106], Harray[75][106], Harray[76][106], Harray[77][106], Harray[78][106], Harray[79][106], Harray[80][106], Harray[81][106], Harray[82][106], Harray[83][106], Harray[84][106], Harray[85][106], Harray[86][106], Harray[87][106], Harray[88][106], Harray[89][106], Harray[90][106], Harray[91][106], Harray[92][106], Harray[93][106], Harray[94][106], Harray[95][106], Harray[96][106], Harray[97][106], Harray[98][106], Harray[99][106], Harray[100][106], Harray[101][106], Harray[102][106], Harray[103][106], Harray[104][106], Harray[105][106], Harray[106][106], Harray[107][106], Harray[108][106], Harray[109][106], Harray[110][106], Harray[111][106], Harray[112][106], Harray[113][106], Harray[114][106], Harray[115][106], Harray[116][106], Harray[117][106], Harray[118][106], Harray[119][106], Harray[120][106], Harray[121][106], Harray[122][106], Harray[123][106], Harray[124][106], Harray[125][106], Harray[126][106], Harray[127][106]};
assign h_col_107 = {Harray[0][107], Harray[1][107], Harray[2][107], Harray[3][107], Harray[4][107], Harray[5][107], Harray[6][107], Harray[7][107], Harray[8][107], Harray[9][107], Harray[10][107], Harray[11][107], Harray[12][107], Harray[13][107], Harray[14][107], Harray[15][107], Harray[16][107], Harray[17][107], Harray[18][107], Harray[19][107], Harray[20][107], Harray[21][107], Harray[22][107], Harray[23][107], Harray[24][107], Harray[25][107], Harray[26][107], Harray[27][107], Harray[28][107], Harray[29][107], Harray[30][107], Harray[31][107], Harray[32][107], Harray[33][107], Harray[34][107], Harray[35][107], Harray[36][107], Harray[37][107], Harray[38][107], Harray[39][107], Harray[40][107], Harray[41][107], Harray[42][107], Harray[43][107], Harray[44][107], Harray[45][107], Harray[46][107], Harray[47][107], Harray[48][107], Harray[49][107], Harray[50][107], Harray[51][107], Harray[52][107], Harray[53][107], Harray[54][107], Harray[55][107], Harray[56][107], Harray[57][107], Harray[58][107], Harray[59][107], Harray[60][107], Harray[61][107], Harray[62][107], Harray[63][107], Harray[64][107], Harray[65][107], Harray[66][107], Harray[67][107], Harray[68][107], Harray[69][107], Harray[70][107], Harray[71][107], Harray[72][107], Harray[73][107], Harray[74][107], Harray[75][107], Harray[76][107], Harray[77][107], Harray[78][107], Harray[79][107], Harray[80][107], Harray[81][107], Harray[82][107], Harray[83][107], Harray[84][107], Harray[85][107], Harray[86][107], Harray[87][107], Harray[88][107], Harray[89][107], Harray[90][107], Harray[91][107], Harray[92][107], Harray[93][107], Harray[94][107], Harray[95][107], Harray[96][107], Harray[97][107], Harray[98][107], Harray[99][107], Harray[100][107], Harray[101][107], Harray[102][107], Harray[103][107], Harray[104][107], Harray[105][107], Harray[106][107], Harray[107][107], Harray[108][107], Harray[109][107], Harray[110][107], Harray[111][107], Harray[112][107], Harray[113][107], Harray[114][107], Harray[115][107], Harray[116][107], Harray[117][107], Harray[118][107], Harray[119][107], Harray[120][107], Harray[121][107], Harray[122][107], Harray[123][107], Harray[124][107], Harray[125][107], Harray[126][107], Harray[127][107]};
assign h_col_108 = {Harray[0][108], Harray[1][108], Harray[2][108], Harray[3][108], Harray[4][108], Harray[5][108], Harray[6][108], Harray[7][108], Harray[8][108], Harray[9][108], Harray[10][108], Harray[11][108], Harray[12][108], Harray[13][108], Harray[14][108], Harray[15][108], Harray[16][108], Harray[17][108], Harray[18][108], Harray[19][108], Harray[20][108], Harray[21][108], Harray[22][108], Harray[23][108], Harray[24][108], Harray[25][108], Harray[26][108], Harray[27][108], Harray[28][108], Harray[29][108], Harray[30][108], Harray[31][108], Harray[32][108], Harray[33][108], Harray[34][108], Harray[35][108], Harray[36][108], Harray[37][108], Harray[38][108], Harray[39][108], Harray[40][108], Harray[41][108], Harray[42][108], Harray[43][108], Harray[44][108], Harray[45][108], Harray[46][108], Harray[47][108], Harray[48][108], Harray[49][108], Harray[50][108], Harray[51][108], Harray[52][108], Harray[53][108], Harray[54][108], Harray[55][108], Harray[56][108], Harray[57][108], Harray[58][108], Harray[59][108], Harray[60][108], Harray[61][108], Harray[62][108], Harray[63][108], Harray[64][108], Harray[65][108], Harray[66][108], Harray[67][108], Harray[68][108], Harray[69][108], Harray[70][108], Harray[71][108], Harray[72][108], Harray[73][108], Harray[74][108], Harray[75][108], Harray[76][108], Harray[77][108], Harray[78][108], Harray[79][108], Harray[80][108], Harray[81][108], Harray[82][108], Harray[83][108], Harray[84][108], Harray[85][108], Harray[86][108], Harray[87][108], Harray[88][108], Harray[89][108], Harray[90][108], Harray[91][108], Harray[92][108], Harray[93][108], Harray[94][108], Harray[95][108], Harray[96][108], Harray[97][108], Harray[98][108], Harray[99][108], Harray[100][108], Harray[101][108], Harray[102][108], Harray[103][108], Harray[104][108], Harray[105][108], Harray[106][108], Harray[107][108], Harray[108][108], Harray[109][108], Harray[110][108], Harray[111][108], Harray[112][108], Harray[113][108], Harray[114][108], Harray[115][108], Harray[116][108], Harray[117][108], Harray[118][108], Harray[119][108], Harray[120][108], Harray[121][108], Harray[122][108], Harray[123][108], Harray[124][108], Harray[125][108], Harray[126][108], Harray[127][108]};
assign h_col_109 = {Harray[0][109], Harray[1][109], Harray[2][109], Harray[3][109], Harray[4][109], Harray[5][109], Harray[6][109], Harray[7][109], Harray[8][109], Harray[9][109], Harray[10][109], Harray[11][109], Harray[12][109], Harray[13][109], Harray[14][109], Harray[15][109], Harray[16][109], Harray[17][109], Harray[18][109], Harray[19][109], Harray[20][109], Harray[21][109], Harray[22][109], Harray[23][109], Harray[24][109], Harray[25][109], Harray[26][109], Harray[27][109], Harray[28][109], Harray[29][109], Harray[30][109], Harray[31][109], Harray[32][109], Harray[33][109], Harray[34][109], Harray[35][109], Harray[36][109], Harray[37][109], Harray[38][109], Harray[39][109], Harray[40][109], Harray[41][109], Harray[42][109], Harray[43][109], Harray[44][109], Harray[45][109], Harray[46][109], Harray[47][109], Harray[48][109], Harray[49][109], Harray[50][109], Harray[51][109], Harray[52][109], Harray[53][109], Harray[54][109], Harray[55][109], Harray[56][109], Harray[57][109], Harray[58][109], Harray[59][109], Harray[60][109], Harray[61][109], Harray[62][109], Harray[63][109], Harray[64][109], Harray[65][109], Harray[66][109], Harray[67][109], Harray[68][109], Harray[69][109], Harray[70][109], Harray[71][109], Harray[72][109], Harray[73][109], Harray[74][109], Harray[75][109], Harray[76][109], Harray[77][109], Harray[78][109], Harray[79][109], Harray[80][109], Harray[81][109], Harray[82][109], Harray[83][109], Harray[84][109], Harray[85][109], Harray[86][109], Harray[87][109], Harray[88][109], Harray[89][109], Harray[90][109], Harray[91][109], Harray[92][109], Harray[93][109], Harray[94][109], Harray[95][109], Harray[96][109], Harray[97][109], Harray[98][109], Harray[99][109], Harray[100][109], Harray[101][109], Harray[102][109], Harray[103][109], Harray[104][109], Harray[105][109], Harray[106][109], Harray[107][109], Harray[108][109], Harray[109][109], Harray[110][109], Harray[111][109], Harray[112][109], Harray[113][109], Harray[114][109], Harray[115][109], Harray[116][109], Harray[117][109], Harray[118][109], Harray[119][109], Harray[120][109], Harray[121][109], Harray[122][109], Harray[123][109], Harray[124][109], Harray[125][109], Harray[126][109], Harray[127][109]};
assign h_col_110 = {Harray[0][110], Harray[1][110], Harray[2][110], Harray[3][110], Harray[4][110], Harray[5][110], Harray[6][110], Harray[7][110], Harray[8][110], Harray[9][110], Harray[10][110], Harray[11][110], Harray[12][110], Harray[13][110], Harray[14][110], Harray[15][110], Harray[16][110], Harray[17][110], Harray[18][110], Harray[19][110], Harray[20][110], Harray[21][110], Harray[22][110], Harray[23][110], Harray[24][110], Harray[25][110], Harray[26][110], Harray[27][110], Harray[28][110], Harray[29][110], Harray[30][110], Harray[31][110], Harray[32][110], Harray[33][110], Harray[34][110], Harray[35][110], Harray[36][110], Harray[37][110], Harray[38][110], Harray[39][110], Harray[40][110], Harray[41][110], Harray[42][110], Harray[43][110], Harray[44][110], Harray[45][110], Harray[46][110], Harray[47][110], Harray[48][110], Harray[49][110], Harray[50][110], Harray[51][110], Harray[52][110], Harray[53][110], Harray[54][110], Harray[55][110], Harray[56][110], Harray[57][110], Harray[58][110], Harray[59][110], Harray[60][110], Harray[61][110], Harray[62][110], Harray[63][110], Harray[64][110], Harray[65][110], Harray[66][110], Harray[67][110], Harray[68][110], Harray[69][110], Harray[70][110], Harray[71][110], Harray[72][110], Harray[73][110], Harray[74][110], Harray[75][110], Harray[76][110], Harray[77][110], Harray[78][110], Harray[79][110], Harray[80][110], Harray[81][110], Harray[82][110], Harray[83][110], Harray[84][110], Harray[85][110], Harray[86][110], Harray[87][110], Harray[88][110], Harray[89][110], Harray[90][110], Harray[91][110], Harray[92][110], Harray[93][110], Harray[94][110], Harray[95][110], Harray[96][110], Harray[97][110], Harray[98][110], Harray[99][110], Harray[100][110], Harray[101][110], Harray[102][110], Harray[103][110], Harray[104][110], Harray[105][110], Harray[106][110], Harray[107][110], Harray[108][110], Harray[109][110], Harray[110][110], Harray[111][110], Harray[112][110], Harray[113][110], Harray[114][110], Harray[115][110], Harray[116][110], Harray[117][110], Harray[118][110], Harray[119][110], Harray[120][110], Harray[121][110], Harray[122][110], Harray[123][110], Harray[124][110], Harray[125][110], Harray[126][110], Harray[127][110]};
assign h_col_111 = {Harray[0][111], Harray[1][111], Harray[2][111], Harray[3][111], Harray[4][111], Harray[5][111], Harray[6][111], Harray[7][111], Harray[8][111], Harray[9][111], Harray[10][111], Harray[11][111], Harray[12][111], Harray[13][111], Harray[14][111], Harray[15][111], Harray[16][111], Harray[17][111], Harray[18][111], Harray[19][111], Harray[20][111], Harray[21][111], Harray[22][111], Harray[23][111], Harray[24][111], Harray[25][111], Harray[26][111], Harray[27][111], Harray[28][111], Harray[29][111], Harray[30][111], Harray[31][111], Harray[32][111], Harray[33][111], Harray[34][111], Harray[35][111], Harray[36][111], Harray[37][111], Harray[38][111], Harray[39][111], Harray[40][111], Harray[41][111], Harray[42][111], Harray[43][111], Harray[44][111], Harray[45][111], Harray[46][111], Harray[47][111], Harray[48][111], Harray[49][111], Harray[50][111], Harray[51][111], Harray[52][111], Harray[53][111], Harray[54][111], Harray[55][111], Harray[56][111], Harray[57][111], Harray[58][111], Harray[59][111], Harray[60][111], Harray[61][111], Harray[62][111], Harray[63][111], Harray[64][111], Harray[65][111], Harray[66][111], Harray[67][111], Harray[68][111], Harray[69][111], Harray[70][111], Harray[71][111], Harray[72][111], Harray[73][111], Harray[74][111], Harray[75][111], Harray[76][111], Harray[77][111], Harray[78][111], Harray[79][111], Harray[80][111], Harray[81][111], Harray[82][111], Harray[83][111], Harray[84][111], Harray[85][111], Harray[86][111], Harray[87][111], Harray[88][111], Harray[89][111], Harray[90][111], Harray[91][111], Harray[92][111], Harray[93][111], Harray[94][111], Harray[95][111], Harray[96][111], Harray[97][111], Harray[98][111], Harray[99][111], Harray[100][111], Harray[101][111], Harray[102][111], Harray[103][111], Harray[104][111], Harray[105][111], Harray[106][111], Harray[107][111], Harray[108][111], Harray[109][111], Harray[110][111], Harray[111][111], Harray[112][111], Harray[113][111], Harray[114][111], Harray[115][111], Harray[116][111], Harray[117][111], Harray[118][111], Harray[119][111], Harray[120][111], Harray[121][111], Harray[122][111], Harray[123][111], Harray[124][111], Harray[125][111], Harray[126][111], Harray[127][111]};
assign h_col_112 = {Harray[0][112], Harray[1][112], Harray[2][112], Harray[3][112], Harray[4][112], Harray[5][112], Harray[6][112], Harray[7][112], Harray[8][112], Harray[9][112], Harray[10][112], Harray[11][112], Harray[12][112], Harray[13][112], Harray[14][112], Harray[15][112], Harray[16][112], Harray[17][112], Harray[18][112], Harray[19][112], Harray[20][112], Harray[21][112], Harray[22][112], Harray[23][112], Harray[24][112], Harray[25][112], Harray[26][112], Harray[27][112], Harray[28][112], Harray[29][112], Harray[30][112], Harray[31][112], Harray[32][112], Harray[33][112], Harray[34][112], Harray[35][112], Harray[36][112], Harray[37][112], Harray[38][112], Harray[39][112], Harray[40][112], Harray[41][112], Harray[42][112], Harray[43][112], Harray[44][112], Harray[45][112], Harray[46][112], Harray[47][112], Harray[48][112], Harray[49][112], Harray[50][112], Harray[51][112], Harray[52][112], Harray[53][112], Harray[54][112], Harray[55][112], Harray[56][112], Harray[57][112], Harray[58][112], Harray[59][112], Harray[60][112], Harray[61][112], Harray[62][112], Harray[63][112], Harray[64][112], Harray[65][112], Harray[66][112], Harray[67][112], Harray[68][112], Harray[69][112], Harray[70][112], Harray[71][112], Harray[72][112], Harray[73][112], Harray[74][112], Harray[75][112], Harray[76][112], Harray[77][112], Harray[78][112], Harray[79][112], Harray[80][112], Harray[81][112], Harray[82][112], Harray[83][112], Harray[84][112], Harray[85][112], Harray[86][112], Harray[87][112], Harray[88][112], Harray[89][112], Harray[90][112], Harray[91][112], Harray[92][112], Harray[93][112], Harray[94][112], Harray[95][112], Harray[96][112], Harray[97][112], Harray[98][112], Harray[99][112], Harray[100][112], Harray[101][112], Harray[102][112], Harray[103][112], Harray[104][112], Harray[105][112], Harray[106][112], Harray[107][112], Harray[108][112], Harray[109][112], Harray[110][112], Harray[111][112], Harray[112][112], Harray[113][112], Harray[114][112], Harray[115][112], Harray[116][112], Harray[117][112], Harray[118][112], Harray[119][112], Harray[120][112], Harray[121][112], Harray[122][112], Harray[123][112], Harray[124][112], Harray[125][112], Harray[126][112], Harray[127][112]};
assign h_col_113 = {Harray[0][113], Harray[1][113], Harray[2][113], Harray[3][113], Harray[4][113], Harray[5][113], Harray[6][113], Harray[7][113], Harray[8][113], Harray[9][113], Harray[10][113], Harray[11][113], Harray[12][113], Harray[13][113], Harray[14][113], Harray[15][113], Harray[16][113], Harray[17][113], Harray[18][113], Harray[19][113], Harray[20][113], Harray[21][113], Harray[22][113], Harray[23][113], Harray[24][113], Harray[25][113], Harray[26][113], Harray[27][113], Harray[28][113], Harray[29][113], Harray[30][113], Harray[31][113], Harray[32][113], Harray[33][113], Harray[34][113], Harray[35][113], Harray[36][113], Harray[37][113], Harray[38][113], Harray[39][113], Harray[40][113], Harray[41][113], Harray[42][113], Harray[43][113], Harray[44][113], Harray[45][113], Harray[46][113], Harray[47][113], Harray[48][113], Harray[49][113], Harray[50][113], Harray[51][113], Harray[52][113], Harray[53][113], Harray[54][113], Harray[55][113], Harray[56][113], Harray[57][113], Harray[58][113], Harray[59][113], Harray[60][113], Harray[61][113], Harray[62][113], Harray[63][113], Harray[64][113], Harray[65][113], Harray[66][113], Harray[67][113], Harray[68][113], Harray[69][113], Harray[70][113], Harray[71][113], Harray[72][113], Harray[73][113], Harray[74][113], Harray[75][113], Harray[76][113], Harray[77][113], Harray[78][113], Harray[79][113], Harray[80][113], Harray[81][113], Harray[82][113], Harray[83][113], Harray[84][113], Harray[85][113], Harray[86][113], Harray[87][113], Harray[88][113], Harray[89][113], Harray[90][113], Harray[91][113], Harray[92][113], Harray[93][113], Harray[94][113], Harray[95][113], Harray[96][113], Harray[97][113], Harray[98][113], Harray[99][113], Harray[100][113], Harray[101][113], Harray[102][113], Harray[103][113], Harray[104][113], Harray[105][113], Harray[106][113], Harray[107][113], Harray[108][113], Harray[109][113], Harray[110][113], Harray[111][113], Harray[112][113], Harray[113][113], Harray[114][113], Harray[115][113], Harray[116][113], Harray[117][113], Harray[118][113], Harray[119][113], Harray[120][113], Harray[121][113], Harray[122][113], Harray[123][113], Harray[124][113], Harray[125][113], Harray[126][113], Harray[127][113]};
assign h_col_114 = {Harray[0][114], Harray[1][114], Harray[2][114], Harray[3][114], Harray[4][114], Harray[5][114], Harray[6][114], Harray[7][114], Harray[8][114], Harray[9][114], Harray[10][114], Harray[11][114], Harray[12][114], Harray[13][114], Harray[14][114], Harray[15][114], Harray[16][114], Harray[17][114], Harray[18][114], Harray[19][114], Harray[20][114], Harray[21][114], Harray[22][114], Harray[23][114], Harray[24][114], Harray[25][114], Harray[26][114], Harray[27][114], Harray[28][114], Harray[29][114], Harray[30][114], Harray[31][114], Harray[32][114], Harray[33][114], Harray[34][114], Harray[35][114], Harray[36][114], Harray[37][114], Harray[38][114], Harray[39][114], Harray[40][114], Harray[41][114], Harray[42][114], Harray[43][114], Harray[44][114], Harray[45][114], Harray[46][114], Harray[47][114], Harray[48][114], Harray[49][114], Harray[50][114], Harray[51][114], Harray[52][114], Harray[53][114], Harray[54][114], Harray[55][114], Harray[56][114], Harray[57][114], Harray[58][114], Harray[59][114], Harray[60][114], Harray[61][114], Harray[62][114], Harray[63][114], Harray[64][114], Harray[65][114], Harray[66][114], Harray[67][114], Harray[68][114], Harray[69][114], Harray[70][114], Harray[71][114], Harray[72][114], Harray[73][114], Harray[74][114], Harray[75][114], Harray[76][114], Harray[77][114], Harray[78][114], Harray[79][114], Harray[80][114], Harray[81][114], Harray[82][114], Harray[83][114], Harray[84][114], Harray[85][114], Harray[86][114], Harray[87][114], Harray[88][114], Harray[89][114], Harray[90][114], Harray[91][114], Harray[92][114], Harray[93][114], Harray[94][114], Harray[95][114], Harray[96][114], Harray[97][114], Harray[98][114], Harray[99][114], Harray[100][114], Harray[101][114], Harray[102][114], Harray[103][114], Harray[104][114], Harray[105][114], Harray[106][114], Harray[107][114], Harray[108][114], Harray[109][114], Harray[110][114], Harray[111][114], Harray[112][114], Harray[113][114], Harray[114][114], Harray[115][114], Harray[116][114], Harray[117][114], Harray[118][114], Harray[119][114], Harray[120][114], Harray[121][114], Harray[122][114], Harray[123][114], Harray[124][114], Harray[125][114], Harray[126][114], Harray[127][114]};
assign h_col_115 = {Harray[0][115], Harray[1][115], Harray[2][115], Harray[3][115], Harray[4][115], Harray[5][115], Harray[6][115], Harray[7][115], Harray[8][115], Harray[9][115], Harray[10][115], Harray[11][115], Harray[12][115], Harray[13][115], Harray[14][115], Harray[15][115], Harray[16][115], Harray[17][115], Harray[18][115], Harray[19][115], Harray[20][115], Harray[21][115], Harray[22][115], Harray[23][115], Harray[24][115], Harray[25][115], Harray[26][115], Harray[27][115], Harray[28][115], Harray[29][115], Harray[30][115], Harray[31][115], Harray[32][115], Harray[33][115], Harray[34][115], Harray[35][115], Harray[36][115], Harray[37][115], Harray[38][115], Harray[39][115], Harray[40][115], Harray[41][115], Harray[42][115], Harray[43][115], Harray[44][115], Harray[45][115], Harray[46][115], Harray[47][115], Harray[48][115], Harray[49][115], Harray[50][115], Harray[51][115], Harray[52][115], Harray[53][115], Harray[54][115], Harray[55][115], Harray[56][115], Harray[57][115], Harray[58][115], Harray[59][115], Harray[60][115], Harray[61][115], Harray[62][115], Harray[63][115], Harray[64][115], Harray[65][115], Harray[66][115], Harray[67][115], Harray[68][115], Harray[69][115], Harray[70][115], Harray[71][115], Harray[72][115], Harray[73][115], Harray[74][115], Harray[75][115], Harray[76][115], Harray[77][115], Harray[78][115], Harray[79][115], Harray[80][115], Harray[81][115], Harray[82][115], Harray[83][115], Harray[84][115], Harray[85][115], Harray[86][115], Harray[87][115], Harray[88][115], Harray[89][115], Harray[90][115], Harray[91][115], Harray[92][115], Harray[93][115], Harray[94][115], Harray[95][115], Harray[96][115], Harray[97][115], Harray[98][115], Harray[99][115], Harray[100][115], Harray[101][115], Harray[102][115], Harray[103][115], Harray[104][115], Harray[105][115], Harray[106][115], Harray[107][115], Harray[108][115], Harray[109][115], Harray[110][115], Harray[111][115], Harray[112][115], Harray[113][115], Harray[114][115], Harray[115][115], Harray[116][115], Harray[117][115], Harray[118][115], Harray[119][115], Harray[120][115], Harray[121][115], Harray[122][115], Harray[123][115], Harray[124][115], Harray[125][115], Harray[126][115], Harray[127][115]};
assign h_col_116 = {Harray[0][116], Harray[1][116], Harray[2][116], Harray[3][116], Harray[4][116], Harray[5][116], Harray[6][116], Harray[7][116], Harray[8][116], Harray[9][116], Harray[10][116], Harray[11][116], Harray[12][116], Harray[13][116], Harray[14][116], Harray[15][116], Harray[16][116], Harray[17][116], Harray[18][116], Harray[19][116], Harray[20][116], Harray[21][116], Harray[22][116], Harray[23][116], Harray[24][116], Harray[25][116], Harray[26][116], Harray[27][116], Harray[28][116], Harray[29][116], Harray[30][116], Harray[31][116], Harray[32][116], Harray[33][116], Harray[34][116], Harray[35][116], Harray[36][116], Harray[37][116], Harray[38][116], Harray[39][116], Harray[40][116], Harray[41][116], Harray[42][116], Harray[43][116], Harray[44][116], Harray[45][116], Harray[46][116], Harray[47][116], Harray[48][116], Harray[49][116], Harray[50][116], Harray[51][116], Harray[52][116], Harray[53][116], Harray[54][116], Harray[55][116], Harray[56][116], Harray[57][116], Harray[58][116], Harray[59][116], Harray[60][116], Harray[61][116], Harray[62][116], Harray[63][116], Harray[64][116], Harray[65][116], Harray[66][116], Harray[67][116], Harray[68][116], Harray[69][116], Harray[70][116], Harray[71][116], Harray[72][116], Harray[73][116], Harray[74][116], Harray[75][116], Harray[76][116], Harray[77][116], Harray[78][116], Harray[79][116], Harray[80][116], Harray[81][116], Harray[82][116], Harray[83][116], Harray[84][116], Harray[85][116], Harray[86][116], Harray[87][116], Harray[88][116], Harray[89][116], Harray[90][116], Harray[91][116], Harray[92][116], Harray[93][116], Harray[94][116], Harray[95][116], Harray[96][116], Harray[97][116], Harray[98][116], Harray[99][116], Harray[100][116], Harray[101][116], Harray[102][116], Harray[103][116], Harray[104][116], Harray[105][116], Harray[106][116], Harray[107][116], Harray[108][116], Harray[109][116], Harray[110][116], Harray[111][116], Harray[112][116], Harray[113][116], Harray[114][116], Harray[115][116], Harray[116][116], Harray[117][116], Harray[118][116], Harray[119][116], Harray[120][116], Harray[121][116], Harray[122][116], Harray[123][116], Harray[124][116], Harray[125][116], Harray[126][116], Harray[127][116]};
assign h_col_117 = {Harray[0][117], Harray[1][117], Harray[2][117], Harray[3][117], Harray[4][117], Harray[5][117], Harray[6][117], Harray[7][117], Harray[8][117], Harray[9][117], Harray[10][117], Harray[11][117], Harray[12][117], Harray[13][117], Harray[14][117], Harray[15][117], Harray[16][117], Harray[17][117], Harray[18][117], Harray[19][117], Harray[20][117], Harray[21][117], Harray[22][117], Harray[23][117], Harray[24][117], Harray[25][117], Harray[26][117], Harray[27][117], Harray[28][117], Harray[29][117], Harray[30][117], Harray[31][117], Harray[32][117], Harray[33][117], Harray[34][117], Harray[35][117], Harray[36][117], Harray[37][117], Harray[38][117], Harray[39][117], Harray[40][117], Harray[41][117], Harray[42][117], Harray[43][117], Harray[44][117], Harray[45][117], Harray[46][117], Harray[47][117], Harray[48][117], Harray[49][117], Harray[50][117], Harray[51][117], Harray[52][117], Harray[53][117], Harray[54][117], Harray[55][117], Harray[56][117], Harray[57][117], Harray[58][117], Harray[59][117], Harray[60][117], Harray[61][117], Harray[62][117], Harray[63][117], Harray[64][117], Harray[65][117], Harray[66][117], Harray[67][117], Harray[68][117], Harray[69][117], Harray[70][117], Harray[71][117], Harray[72][117], Harray[73][117], Harray[74][117], Harray[75][117], Harray[76][117], Harray[77][117], Harray[78][117], Harray[79][117], Harray[80][117], Harray[81][117], Harray[82][117], Harray[83][117], Harray[84][117], Harray[85][117], Harray[86][117], Harray[87][117], Harray[88][117], Harray[89][117], Harray[90][117], Harray[91][117], Harray[92][117], Harray[93][117], Harray[94][117], Harray[95][117], Harray[96][117], Harray[97][117], Harray[98][117], Harray[99][117], Harray[100][117], Harray[101][117], Harray[102][117], Harray[103][117], Harray[104][117], Harray[105][117], Harray[106][117], Harray[107][117], Harray[108][117], Harray[109][117], Harray[110][117], Harray[111][117], Harray[112][117], Harray[113][117], Harray[114][117], Harray[115][117], Harray[116][117], Harray[117][117], Harray[118][117], Harray[119][117], Harray[120][117], Harray[121][117], Harray[122][117], Harray[123][117], Harray[124][117], Harray[125][117], Harray[126][117], Harray[127][117]};
assign h_col_118 = {Harray[0][118], Harray[1][118], Harray[2][118], Harray[3][118], Harray[4][118], Harray[5][118], Harray[6][118], Harray[7][118], Harray[8][118], Harray[9][118], Harray[10][118], Harray[11][118], Harray[12][118], Harray[13][118], Harray[14][118], Harray[15][118], Harray[16][118], Harray[17][118], Harray[18][118], Harray[19][118], Harray[20][118], Harray[21][118], Harray[22][118], Harray[23][118], Harray[24][118], Harray[25][118], Harray[26][118], Harray[27][118], Harray[28][118], Harray[29][118], Harray[30][118], Harray[31][118], Harray[32][118], Harray[33][118], Harray[34][118], Harray[35][118], Harray[36][118], Harray[37][118], Harray[38][118], Harray[39][118], Harray[40][118], Harray[41][118], Harray[42][118], Harray[43][118], Harray[44][118], Harray[45][118], Harray[46][118], Harray[47][118], Harray[48][118], Harray[49][118], Harray[50][118], Harray[51][118], Harray[52][118], Harray[53][118], Harray[54][118], Harray[55][118], Harray[56][118], Harray[57][118], Harray[58][118], Harray[59][118], Harray[60][118], Harray[61][118], Harray[62][118], Harray[63][118], Harray[64][118], Harray[65][118], Harray[66][118], Harray[67][118], Harray[68][118], Harray[69][118], Harray[70][118], Harray[71][118], Harray[72][118], Harray[73][118], Harray[74][118], Harray[75][118], Harray[76][118], Harray[77][118], Harray[78][118], Harray[79][118], Harray[80][118], Harray[81][118], Harray[82][118], Harray[83][118], Harray[84][118], Harray[85][118], Harray[86][118], Harray[87][118], Harray[88][118], Harray[89][118], Harray[90][118], Harray[91][118], Harray[92][118], Harray[93][118], Harray[94][118], Harray[95][118], Harray[96][118], Harray[97][118], Harray[98][118], Harray[99][118], Harray[100][118], Harray[101][118], Harray[102][118], Harray[103][118], Harray[104][118], Harray[105][118], Harray[106][118], Harray[107][118], Harray[108][118], Harray[109][118], Harray[110][118], Harray[111][118], Harray[112][118], Harray[113][118], Harray[114][118], Harray[115][118], Harray[116][118], Harray[117][118], Harray[118][118], Harray[119][118], Harray[120][118], Harray[121][118], Harray[122][118], Harray[123][118], Harray[124][118], Harray[125][118], Harray[126][118], Harray[127][118]};
assign h_col_119 = {Harray[0][119], Harray[1][119], Harray[2][119], Harray[3][119], Harray[4][119], Harray[5][119], Harray[6][119], Harray[7][119], Harray[8][119], Harray[9][119], Harray[10][119], Harray[11][119], Harray[12][119], Harray[13][119], Harray[14][119], Harray[15][119], Harray[16][119], Harray[17][119], Harray[18][119], Harray[19][119], Harray[20][119], Harray[21][119], Harray[22][119], Harray[23][119], Harray[24][119], Harray[25][119], Harray[26][119], Harray[27][119], Harray[28][119], Harray[29][119], Harray[30][119], Harray[31][119], Harray[32][119], Harray[33][119], Harray[34][119], Harray[35][119], Harray[36][119], Harray[37][119], Harray[38][119], Harray[39][119], Harray[40][119], Harray[41][119], Harray[42][119], Harray[43][119], Harray[44][119], Harray[45][119], Harray[46][119], Harray[47][119], Harray[48][119], Harray[49][119], Harray[50][119], Harray[51][119], Harray[52][119], Harray[53][119], Harray[54][119], Harray[55][119], Harray[56][119], Harray[57][119], Harray[58][119], Harray[59][119], Harray[60][119], Harray[61][119], Harray[62][119], Harray[63][119], Harray[64][119], Harray[65][119], Harray[66][119], Harray[67][119], Harray[68][119], Harray[69][119], Harray[70][119], Harray[71][119], Harray[72][119], Harray[73][119], Harray[74][119], Harray[75][119], Harray[76][119], Harray[77][119], Harray[78][119], Harray[79][119], Harray[80][119], Harray[81][119], Harray[82][119], Harray[83][119], Harray[84][119], Harray[85][119], Harray[86][119], Harray[87][119], Harray[88][119], Harray[89][119], Harray[90][119], Harray[91][119], Harray[92][119], Harray[93][119], Harray[94][119], Harray[95][119], Harray[96][119], Harray[97][119], Harray[98][119], Harray[99][119], Harray[100][119], Harray[101][119], Harray[102][119], Harray[103][119], Harray[104][119], Harray[105][119], Harray[106][119], Harray[107][119], Harray[108][119], Harray[109][119], Harray[110][119], Harray[111][119], Harray[112][119], Harray[113][119], Harray[114][119], Harray[115][119], Harray[116][119], Harray[117][119], Harray[118][119], Harray[119][119], Harray[120][119], Harray[121][119], Harray[122][119], Harray[123][119], Harray[124][119], Harray[125][119], Harray[126][119], Harray[127][119]};
assign h_col_120 = {Harray[0][120], Harray[1][120], Harray[2][120], Harray[3][120], Harray[4][120], Harray[5][120], Harray[6][120], Harray[7][120], Harray[8][120], Harray[9][120], Harray[10][120], Harray[11][120], Harray[12][120], Harray[13][120], Harray[14][120], Harray[15][120], Harray[16][120], Harray[17][120], Harray[18][120], Harray[19][120], Harray[20][120], Harray[21][120], Harray[22][120], Harray[23][120], Harray[24][120], Harray[25][120], Harray[26][120], Harray[27][120], Harray[28][120], Harray[29][120], Harray[30][120], Harray[31][120], Harray[32][120], Harray[33][120], Harray[34][120], Harray[35][120], Harray[36][120], Harray[37][120], Harray[38][120], Harray[39][120], Harray[40][120], Harray[41][120], Harray[42][120], Harray[43][120], Harray[44][120], Harray[45][120], Harray[46][120], Harray[47][120], Harray[48][120], Harray[49][120], Harray[50][120], Harray[51][120], Harray[52][120], Harray[53][120], Harray[54][120], Harray[55][120], Harray[56][120], Harray[57][120], Harray[58][120], Harray[59][120], Harray[60][120], Harray[61][120], Harray[62][120], Harray[63][120], Harray[64][120], Harray[65][120], Harray[66][120], Harray[67][120], Harray[68][120], Harray[69][120], Harray[70][120], Harray[71][120], Harray[72][120], Harray[73][120], Harray[74][120], Harray[75][120], Harray[76][120], Harray[77][120], Harray[78][120], Harray[79][120], Harray[80][120], Harray[81][120], Harray[82][120], Harray[83][120], Harray[84][120], Harray[85][120], Harray[86][120], Harray[87][120], Harray[88][120], Harray[89][120], Harray[90][120], Harray[91][120], Harray[92][120], Harray[93][120], Harray[94][120], Harray[95][120], Harray[96][120], Harray[97][120], Harray[98][120], Harray[99][120], Harray[100][120], Harray[101][120], Harray[102][120], Harray[103][120], Harray[104][120], Harray[105][120], Harray[106][120], Harray[107][120], Harray[108][120], Harray[109][120], Harray[110][120], Harray[111][120], Harray[112][120], Harray[113][120], Harray[114][120], Harray[115][120], Harray[116][120], Harray[117][120], Harray[118][120], Harray[119][120], Harray[120][120], Harray[121][120], Harray[122][120], Harray[123][120], Harray[124][120], Harray[125][120], Harray[126][120], Harray[127][120]};
assign h_col_121 = {Harray[0][121], Harray[1][121], Harray[2][121], Harray[3][121], Harray[4][121], Harray[5][121], Harray[6][121], Harray[7][121], Harray[8][121], Harray[9][121], Harray[10][121], Harray[11][121], Harray[12][121], Harray[13][121], Harray[14][121], Harray[15][121], Harray[16][121], Harray[17][121], Harray[18][121], Harray[19][121], Harray[20][121], Harray[21][121], Harray[22][121], Harray[23][121], Harray[24][121], Harray[25][121], Harray[26][121], Harray[27][121], Harray[28][121], Harray[29][121], Harray[30][121], Harray[31][121], Harray[32][121], Harray[33][121], Harray[34][121], Harray[35][121], Harray[36][121], Harray[37][121], Harray[38][121], Harray[39][121], Harray[40][121], Harray[41][121], Harray[42][121], Harray[43][121], Harray[44][121], Harray[45][121], Harray[46][121], Harray[47][121], Harray[48][121], Harray[49][121], Harray[50][121], Harray[51][121], Harray[52][121], Harray[53][121], Harray[54][121], Harray[55][121], Harray[56][121], Harray[57][121], Harray[58][121], Harray[59][121], Harray[60][121], Harray[61][121], Harray[62][121], Harray[63][121], Harray[64][121], Harray[65][121], Harray[66][121], Harray[67][121], Harray[68][121], Harray[69][121], Harray[70][121], Harray[71][121], Harray[72][121], Harray[73][121], Harray[74][121], Harray[75][121], Harray[76][121], Harray[77][121], Harray[78][121], Harray[79][121], Harray[80][121], Harray[81][121], Harray[82][121], Harray[83][121], Harray[84][121], Harray[85][121], Harray[86][121], Harray[87][121], Harray[88][121], Harray[89][121], Harray[90][121], Harray[91][121], Harray[92][121], Harray[93][121], Harray[94][121], Harray[95][121], Harray[96][121], Harray[97][121], Harray[98][121], Harray[99][121], Harray[100][121], Harray[101][121], Harray[102][121], Harray[103][121], Harray[104][121], Harray[105][121], Harray[106][121], Harray[107][121], Harray[108][121], Harray[109][121], Harray[110][121], Harray[111][121], Harray[112][121], Harray[113][121], Harray[114][121], Harray[115][121], Harray[116][121], Harray[117][121], Harray[118][121], Harray[119][121], Harray[120][121], Harray[121][121], Harray[122][121], Harray[123][121], Harray[124][121], Harray[125][121], Harray[126][121], Harray[127][121]};
assign h_col_122 = {Harray[0][122], Harray[1][122], Harray[2][122], Harray[3][122], Harray[4][122], Harray[5][122], Harray[6][122], Harray[7][122], Harray[8][122], Harray[9][122], Harray[10][122], Harray[11][122], Harray[12][122], Harray[13][122], Harray[14][122], Harray[15][122], Harray[16][122], Harray[17][122], Harray[18][122], Harray[19][122], Harray[20][122], Harray[21][122], Harray[22][122], Harray[23][122], Harray[24][122], Harray[25][122], Harray[26][122], Harray[27][122], Harray[28][122], Harray[29][122], Harray[30][122], Harray[31][122], Harray[32][122], Harray[33][122], Harray[34][122], Harray[35][122], Harray[36][122], Harray[37][122], Harray[38][122], Harray[39][122], Harray[40][122], Harray[41][122], Harray[42][122], Harray[43][122], Harray[44][122], Harray[45][122], Harray[46][122], Harray[47][122], Harray[48][122], Harray[49][122], Harray[50][122], Harray[51][122], Harray[52][122], Harray[53][122], Harray[54][122], Harray[55][122], Harray[56][122], Harray[57][122], Harray[58][122], Harray[59][122], Harray[60][122], Harray[61][122], Harray[62][122], Harray[63][122], Harray[64][122], Harray[65][122], Harray[66][122], Harray[67][122], Harray[68][122], Harray[69][122], Harray[70][122], Harray[71][122], Harray[72][122], Harray[73][122], Harray[74][122], Harray[75][122], Harray[76][122], Harray[77][122], Harray[78][122], Harray[79][122], Harray[80][122], Harray[81][122], Harray[82][122], Harray[83][122], Harray[84][122], Harray[85][122], Harray[86][122], Harray[87][122], Harray[88][122], Harray[89][122], Harray[90][122], Harray[91][122], Harray[92][122], Harray[93][122], Harray[94][122], Harray[95][122], Harray[96][122], Harray[97][122], Harray[98][122], Harray[99][122], Harray[100][122], Harray[101][122], Harray[102][122], Harray[103][122], Harray[104][122], Harray[105][122], Harray[106][122], Harray[107][122], Harray[108][122], Harray[109][122], Harray[110][122], Harray[111][122], Harray[112][122], Harray[113][122], Harray[114][122], Harray[115][122], Harray[116][122], Harray[117][122], Harray[118][122], Harray[119][122], Harray[120][122], Harray[121][122], Harray[122][122], Harray[123][122], Harray[124][122], Harray[125][122], Harray[126][122], Harray[127][122]};
assign h_col_123 = {Harray[0][123], Harray[1][123], Harray[2][123], Harray[3][123], Harray[4][123], Harray[5][123], Harray[6][123], Harray[7][123], Harray[8][123], Harray[9][123], Harray[10][123], Harray[11][123], Harray[12][123], Harray[13][123], Harray[14][123], Harray[15][123], Harray[16][123], Harray[17][123], Harray[18][123], Harray[19][123], Harray[20][123], Harray[21][123], Harray[22][123], Harray[23][123], Harray[24][123], Harray[25][123], Harray[26][123], Harray[27][123], Harray[28][123], Harray[29][123], Harray[30][123], Harray[31][123], Harray[32][123], Harray[33][123], Harray[34][123], Harray[35][123], Harray[36][123], Harray[37][123], Harray[38][123], Harray[39][123], Harray[40][123], Harray[41][123], Harray[42][123], Harray[43][123], Harray[44][123], Harray[45][123], Harray[46][123], Harray[47][123], Harray[48][123], Harray[49][123], Harray[50][123], Harray[51][123], Harray[52][123], Harray[53][123], Harray[54][123], Harray[55][123], Harray[56][123], Harray[57][123], Harray[58][123], Harray[59][123], Harray[60][123], Harray[61][123], Harray[62][123], Harray[63][123], Harray[64][123], Harray[65][123], Harray[66][123], Harray[67][123], Harray[68][123], Harray[69][123], Harray[70][123], Harray[71][123], Harray[72][123], Harray[73][123], Harray[74][123], Harray[75][123], Harray[76][123], Harray[77][123], Harray[78][123], Harray[79][123], Harray[80][123], Harray[81][123], Harray[82][123], Harray[83][123], Harray[84][123], Harray[85][123], Harray[86][123], Harray[87][123], Harray[88][123], Harray[89][123], Harray[90][123], Harray[91][123], Harray[92][123], Harray[93][123], Harray[94][123], Harray[95][123], Harray[96][123], Harray[97][123], Harray[98][123], Harray[99][123], Harray[100][123], Harray[101][123], Harray[102][123], Harray[103][123], Harray[104][123], Harray[105][123], Harray[106][123], Harray[107][123], Harray[108][123], Harray[109][123], Harray[110][123], Harray[111][123], Harray[112][123], Harray[113][123], Harray[114][123], Harray[115][123], Harray[116][123], Harray[117][123], Harray[118][123], Harray[119][123], Harray[120][123], Harray[121][123], Harray[122][123], Harray[123][123], Harray[124][123], Harray[125][123], Harray[126][123], Harray[127][123]};
assign h_col_124 = {Harray[0][124], Harray[1][124], Harray[2][124], Harray[3][124], Harray[4][124], Harray[5][124], Harray[6][124], Harray[7][124], Harray[8][124], Harray[9][124], Harray[10][124], Harray[11][124], Harray[12][124], Harray[13][124], Harray[14][124], Harray[15][124], Harray[16][124], Harray[17][124], Harray[18][124], Harray[19][124], Harray[20][124], Harray[21][124], Harray[22][124], Harray[23][124], Harray[24][124], Harray[25][124], Harray[26][124], Harray[27][124], Harray[28][124], Harray[29][124], Harray[30][124], Harray[31][124], Harray[32][124], Harray[33][124], Harray[34][124], Harray[35][124], Harray[36][124], Harray[37][124], Harray[38][124], Harray[39][124], Harray[40][124], Harray[41][124], Harray[42][124], Harray[43][124], Harray[44][124], Harray[45][124], Harray[46][124], Harray[47][124], Harray[48][124], Harray[49][124], Harray[50][124], Harray[51][124], Harray[52][124], Harray[53][124], Harray[54][124], Harray[55][124], Harray[56][124], Harray[57][124], Harray[58][124], Harray[59][124], Harray[60][124], Harray[61][124], Harray[62][124], Harray[63][124], Harray[64][124], Harray[65][124], Harray[66][124], Harray[67][124], Harray[68][124], Harray[69][124], Harray[70][124], Harray[71][124], Harray[72][124], Harray[73][124], Harray[74][124], Harray[75][124], Harray[76][124], Harray[77][124], Harray[78][124], Harray[79][124], Harray[80][124], Harray[81][124], Harray[82][124], Harray[83][124], Harray[84][124], Harray[85][124], Harray[86][124], Harray[87][124], Harray[88][124], Harray[89][124], Harray[90][124], Harray[91][124], Harray[92][124], Harray[93][124], Harray[94][124], Harray[95][124], Harray[96][124], Harray[97][124], Harray[98][124], Harray[99][124], Harray[100][124], Harray[101][124], Harray[102][124], Harray[103][124], Harray[104][124], Harray[105][124], Harray[106][124], Harray[107][124], Harray[108][124], Harray[109][124], Harray[110][124], Harray[111][124], Harray[112][124], Harray[113][124], Harray[114][124], Harray[115][124], Harray[116][124], Harray[117][124], Harray[118][124], Harray[119][124], Harray[120][124], Harray[121][124], Harray[122][124], Harray[123][124], Harray[124][124], Harray[125][124], Harray[126][124], Harray[127][124]};
assign h_col_125 = {Harray[0][125], Harray[1][125], Harray[2][125], Harray[3][125], Harray[4][125], Harray[5][125], Harray[6][125], Harray[7][125], Harray[8][125], Harray[9][125], Harray[10][125], Harray[11][125], Harray[12][125], Harray[13][125], Harray[14][125], Harray[15][125], Harray[16][125], Harray[17][125], Harray[18][125], Harray[19][125], Harray[20][125], Harray[21][125], Harray[22][125], Harray[23][125], Harray[24][125], Harray[25][125], Harray[26][125], Harray[27][125], Harray[28][125], Harray[29][125], Harray[30][125], Harray[31][125], Harray[32][125], Harray[33][125], Harray[34][125], Harray[35][125], Harray[36][125], Harray[37][125], Harray[38][125], Harray[39][125], Harray[40][125], Harray[41][125], Harray[42][125], Harray[43][125], Harray[44][125], Harray[45][125], Harray[46][125], Harray[47][125], Harray[48][125], Harray[49][125], Harray[50][125], Harray[51][125], Harray[52][125], Harray[53][125], Harray[54][125], Harray[55][125], Harray[56][125], Harray[57][125], Harray[58][125], Harray[59][125], Harray[60][125], Harray[61][125], Harray[62][125], Harray[63][125], Harray[64][125], Harray[65][125], Harray[66][125], Harray[67][125], Harray[68][125], Harray[69][125], Harray[70][125], Harray[71][125], Harray[72][125], Harray[73][125], Harray[74][125], Harray[75][125], Harray[76][125], Harray[77][125], Harray[78][125], Harray[79][125], Harray[80][125], Harray[81][125], Harray[82][125], Harray[83][125], Harray[84][125], Harray[85][125], Harray[86][125], Harray[87][125], Harray[88][125], Harray[89][125], Harray[90][125], Harray[91][125], Harray[92][125], Harray[93][125], Harray[94][125], Harray[95][125], Harray[96][125], Harray[97][125], Harray[98][125], Harray[99][125], Harray[100][125], Harray[101][125], Harray[102][125], Harray[103][125], Harray[104][125], Harray[105][125], Harray[106][125], Harray[107][125], Harray[108][125], Harray[109][125], Harray[110][125], Harray[111][125], Harray[112][125], Harray[113][125], Harray[114][125], Harray[115][125], Harray[116][125], Harray[117][125], Harray[118][125], Harray[119][125], Harray[120][125], Harray[121][125], Harray[122][125], Harray[123][125], Harray[124][125], Harray[125][125], Harray[126][125], Harray[127][125]};
assign h_col_126 = {Harray[0][126], Harray[1][126], Harray[2][126], Harray[3][126], Harray[4][126], Harray[5][126], Harray[6][126], Harray[7][126], Harray[8][126], Harray[9][126], Harray[10][126], Harray[11][126], Harray[12][126], Harray[13][126], Harray[14][126], Harray[15][126], Harray[16][126], Harray[17][126], Harray[18][126], Harray[19][126], Harray[20][126], Harray[21][126], Harray[22][126], Harray[23][126], Harray[24][126], Harray[25][126], Harray[26][126], Harray[27][126], Harray[28][126], Harray[29][126], Harray[30][126], Harray[31][126], Harray[32][126], Harray[33][126], Harray[34][126], Harray[35][126], Harray[36][126], Harray[37][126], Harray[38][126], Harray[39][126], Harray[40][126], Harray[41][126], Harray[42][126], Harray[43][126], Harray[44][126], Harray[45][126], Harray[46][126], Harray[47][126], Harray[48][126], Harray[49][126], Harray[50][126], Harray[51][126], Harray[52][126], Harray[53][126], Harray[54][126], Harray[55][126], Harray[56][126], Harray[57][126], Harray[58][126], Harray[59][126], Harray[60][126], Harray[61][126], Harray[62][126], Harray[63][126], Harray[64][126], Harray[65][126], Harray[66][126], Harray[67][126], Harray[68][126], Harray[69][126], Harray[70][126], Harray[71][126], Harray[72][126], Harray[73][126], Harray[74][126], Harray[75][126], Harray[76][126], Harray[77][126], Harray[78][126], Harray[79][126], Harray[80][126], Harray[81][126], Harray[82][126], Harray[83][126], Harray[84][126], Harray[85][126], Harray[86][126], Harray[87][126], Harray[88][126], Harray[89][126], Harray[90][126], Harray[91][126], Harray[92][126], Harray[93][126], Harray[94][126], Harray[95][126], Harray[96][126], Harray[97][126], Harray[98][126], Harray[99][126], Harray[100][126], Harray[101][126], Harray[102][126], Harray[103][126], Harray[104][126], Harray[105][126], Harray[106][126], Harray[107][126], Harray[108][126], Harray[109][126], Harray[110][126], Harray[111][126], Harray[112][126], Harray[113][126], Harray[114][126], Harray[115][126], Harray[116][126], Harray[117][126], Harray[118][126], Harray[119][126], Harray[120][126], Harray[121][126], Harray[122][126], Harray[123][126], Harray[124][126], Harray[125][126], Harray[126][126], Harray[127][126]};
assign h_col_127 = {Harray[0][127], Harray[1][127], Harray[2][127], Harray[3][127], Harray[4][127], Harray[5][127], Harray[6][127], Harray[7][127], Harray[8][127], Harray[9][127], Harray[10][127], Harray[11][127], Harray[12][127], Harray[13][127], Harray[14][127], Harray[15][127], Harray[16][127], Harray[17][127], Harray[18][127], Harray[19][127], Harray[20][127], Harray[21][127], Harray[22][127], Harray[23][127], Harray[24][127], Harray[25][127], Harray[26][127], Harray[27][127], Harray[28][127], Harray[29][127], Harray[30][127], Harray[31][127], Harray[32][127], Harray[33][127], Harray[34][127], Harray[35][127], Harray[36][127], Harray[37][127], Harray[38][127], Harray[39][127], Harray[40][127], Harray[41][127], Harray[42][127], Harray[43][127], Harray[44][127], Harray[45][127], Harray[46][127], Harray[47][127], Harray[48][127], Harray[49][127], Harray[50][127], Harray[51][127], Harray[52][127], Harray[53][127], Harray[54][127], Harray[55][127], Harray[56][127], Harray[57][127], Harray[58][127], Harray[59][127], Harray[60][127], Harray[61][127], Harray[62][127], Harray[63][127], Harray[64][127], Harray[65][127], Harray[66][127], Harray[67][127], Harray[68][127], Harray[69][127], Harray[70][127], Harray[71][127], Harray[72][127], Harray[73][127], Harray[74][127], Harray[75][127], Harray[76][127], Harray[77][127], Harray[78][127], Harray[79][127], Harray[80][127], Harray[81][127], Harray[82][127], Harray[83][127], Harray[84][127], Harray[85][127], Harray[86][127], Harray[87][127], Harray[88][127], Harray[89][127], Harray[90][127], Harray[91][127], Harray[92][127], Harray[93][127], Harray[94][127], Harray[95][127], Harray[96][127], Harray[97][127], Harray[98][127], Harray[99][127], Harray[100][127], Harray[101][127], Harray[102][127], Harray[103][127], Harray[104][127], Harray[105][127], Harray[106][127], Harray[107][127], Harray[108][127], Harray[109][127], Harray[110][127], Harray[111][127], Harray[112][127], Harray[113][127], Harray[114][127], Harray[115][127], Harray[116][127], Harray[117][127], Harray[118][127], Harray[119][127], Harray[120][127], Harray[121][127], Harray[122][127], Harray[123][127], Harray[124][127], Harray[125][127], Harray[126][127], Harray[127][127]};
assign h_col_128 = {Harray[0][128], Harray[1][128], Harray[2][128], Harray[3][128], Harray[4][128], Harray[5][128], Harray[6][128], Harray[7][128], Harray[8][128], Harray[9][128], Harray[10][128], Harray[11][128], Harray[12][128], Harray[13][128], Harray[14][128], Harray[15][128], Harray[16][128], Harray[17][128], Harray[18][128], Harray[19][128], Harray[20][128], Harray[21][128], Harray[22][128], Harray[23][128], Harray[24][128], Harray[25][128], Harray[26][128], Harray[27][128], Harray[28][128], Harray[29][128], Harray[30][128], Harray[31][128], Harray[32][128], Harray[33][128], Harray[34][128], Harray[35][128], Harray[36][128], Harray[37][128], Harray[38][128], Harray[39][128], Harray[40][128], Harray[41][128], Harray[42][128], Harray[43][128], Harray[44][128], Harray[45][128], Harray[46][128], Harray[47][128], Harray[48][128], Harray[49][128], Harray[50][128], Harray[51][128], Harray[52][128], Harray[53][128], Harray[54][128], Harray[55][128], Harray[56][128], Harray[57][128], Harray[58][128], Harray[59][128], Harray[60][128], Harray[61][128], Harray[62][128], Harray[63][128], Harray[64][128], Harray[65][128], Harray[66][128], Harray[67][128], Harray[68][128], Harray[69][128], Harray[70][128], Harray[71][128], Harray[72][128], Harray[73][128], Harray[74][128], Harray[75][128], Harray[76][128], Harray[77][128], Harray[78][128], Harray[79][128], Harray[80][128], Harray[81][128], Harray[82][128], Harray[83][128], Harray[84][128], Harray[85][128], Harray[86][128], Harray[87][128], Harray[88][128], Harray[89][128], Harray[90][128], Harray[91][128], Harray[92][128], Harray[93][128], Harray[94][128], Harray[95][128], Harray[96][128], Harray[97][128], Harray[98][128], Harray[99][128], Harray[100][128], Harray[101][128], Harray[102][128], Harray[103][128], Harray[104][128], Harray[105][128], Harray[106][128], Harray[107][128], Harray[108][128], Harray[109][128], Harray[110][128], Harray[111][128], Harray[112][128], Harray[113][128], Harray[114][128], Harray[115][128], Harray[116][128], Harray[117][128], Harray[118][128], Harray[119][128], Harray[120][128], Harray[121][128], Harray[122][128], Harray[123][128], Harray[124][128], Harray[125][128], Harray[126][128], Harray[127][128]};
assign h_col_129 = {Harray[0][129], Harray[1][129], Harray[2][129], Harray[3][129], Harray[4][129], Harray[5][129], Harray[6][129], Harray[7][129], Harray[8][129], Harray[9][129], Harray[10][129], Harray[11][129], Harray[12][129], Harray[13][129], Harray[14][129], Harray[15][129], Harray[16][129], Harray[17][129], Harray[18][129], Harray[19][129], Harray[20][129], Harray[21][129], Harray[22][129], Harray[23][129], Harray[24][129], Harray[25][129], Harray[26][129], Harray[27][129], Harray[28][129], Harray[29][129], Harray[30][129], Harray[31][129], Harray[32][129], Harray[33][129], Harray[34][129], Harray[35][129], Harray[36][129], Harray[37][129], Harray[38][129], Harray[39][129], Harray[40][129], Harray[41][129], Harray[42][129], Harray[43][129], Harray[44][129], Harray[45][129], Harray[46][129], Harray[47][129], Harray[48][129], Harray[49][129], Harray[50][129], Harray[51][129], Harray[52][129], Harray[53][129], Harray[54][129], Harray[55][129], Harray[56][129], Harray[57][129], Harray[58][129], Harray[59][129], Harray[60][129], Harray[61][129], Harray[62][129], Harray[63][129], Harray[64][129], Harray[65][129], Harray[66][129], Harray[67][129], Harray[68][129], Harray[69][129], Harray[70][129], Harray[71][129], Harray[72][129], Harray[73][129], Harray[74][129], Harray[75][129], Harray[76][129], Harray[77][129], Harray[78][129], Harray[79][129], Harray[80][129], Harray[81][129], Harray[82][129], Harray[83][129], Harray[84][129], Harray[85][129], Harray[86][129], Harray[87][129], Harray[88][129], Harray[89][129], Harray[90][129], Harray[91][129], Harray[92][129], Harray[93][129], Harray[94][129], Harray[95][129], Harray[96][129], Harray[97][129], Harray[98][129], Harray[99][129], Harray[100][129], Harray[101][129], Harray[102][129], Harray[103][129], Harray[104][129], Harray[105][129], Harray[106][129], Harray[107][129], Harray[108][129], Harray[109][129], Harray[110][129], Harray[111][129], Harray[112][129], Harray[113][129], Harray[114][129], Harray[115][129], Harray[116][129], Harray[117][129], Harray[118][129], Harray[119][129], Harray[120][129], Harray[121][129], Harray[122][129], Harray[123][129], Harray[124][129], Harray[125][129], Harray[126][129], Harray[127][129]};
assign h_col_130 = {Harray[0][130], Harray[1][130], Harray[2][130], Harray[3][130], Harray[4][130], Harray[5][130], Harray[6][130], Harray[7][130], Harray[8][130], Harray[9][130], Harray[10][130], Harray[11][130], Harray[12][130], Harray[13][130], Harray[14][130], Harray[15][130], Harray[16][130], Harray[17][130], Harray[18][130], Harray[19][130], Harray[20][130], Harray[21][130], Harray[22][130], Harray[23][130], Harray[24][130], Harray[25][130], Harray[26][130], Harray[27][130], Harray[28][130], Harray[29][130], Harray[30][130], Harray[31][130], Harray[32][130], Harray[33][130], Harray[34][130], Harray[35][130], Harray[36][130], Harray[37][130], Harray[38][130], Harray[39][130], Harray[40][130], Harray[41][130], Harray[42][130], Harray[43][130], Harray[44][130], Harray[45][130], Harray[46][130], Harray[47][130], Harray[48][130], Harray[49][130], Harray[50][130], Harray[51][130], Harray[52][130], Harray[53][130], Harray[54][130], Harray[55][130], Harray[56][130], Harray[57][130], Harray[58][130], Harray[59][130], Harray[60][130], Harray[61][130], Harray[62][130], Harray[63][130], Harray[64][130], Harray[65][130], Harray[66][130], Harray[67][130], Harray[68][130], Harray[69][130], Harray[70][130], Harray[71][130], Harray[72][130], Harray[73][130], Harray[74][130], Harray[75][130], Harray[76][130], Harray[77][130], Harray[78][130], Harray[79][130], Harray[80][130], Harray[81][130], Harray[82][130], Harray[83][130], Harray[84][130], Harray[85][130], Harray[86][130], Harray[87][130], Harray[88][130], Harray[89][130], Harray[90][130], Harray[91][130], Harray[92][130], Harray[93][130], Harray[94][130], Harray[95][130], Harray[96][130], Harray[97][130], Harray[98][130], Harray[99][130], Harray[100][130], Harray[101][130], Harray[102][130], Harray[103][130], Harray[104][130], Harray[105][130], Harray[106][130], Harray[107][130], Harray[108][130], Harray[109][130], Harray[110][130], Harray[111][130], Harray[112][130], Harray[113][130], Harray[114][130], Harray[115][130], Harray[116][130], Harray[117][130], Harray[118][130], Harray[119][130], Harray[120][130], Harray[121][130], Harray[122][130], Harray[123][130], Harray[124][130], Harray[125][130], Harray[126][130], Harray[127][130]};
assign h_col_131 = {Harray[0][131], Harray[1][131], Harray[2][131], Harray[3][131], Harray[4][131], Harray[5][131], Harray[6][131], Harray[7][131], Harray[8][131], Harray[9][131], Harray[10][131], Harray[11][131], Harray[12][131], Harray[13][131], Harray[14][131], Harray[15][131], Harray[16][131], Harray[17][131], Harray[18][131], Harray[19][131], Harray[20][131], Harray[21][131], Harray[22][131], Harray[23][131], Harray[24][131], Harray[25][131], Harray[26][131], Harray[27][131], Harray[28][131], Harray[29][131], Harray[30][131], Harray[31][131], Harray[32][131], Harray[33][131], Harray[34][131], Harray[35][131], Harray[36][131], Harray[37][131], Harray[38][131], Harray[39][131], Harray[40][131], Harray[41][131], Harray[42][131], Harray[43][131], Harray[44][131], Harray[45][131], Harray[46][131], Harray[47][131], Harray[48][131], Harray[49][131], Harray[50][131], Harray[51][131], Harray[52][131], Harray[53][131], Harray[54][131], Harray[55][131], Harray[56][131], Harray[57][131], Harray[58][131], Harray[59][131], Harray[60][131], Harray[61][131], Harray[62][131], Harray[63][131], Harray[64][131], Harray[65][131], Harray[66][131], Harray[67][131], Harray[68][131], Harray[69][131], Harray[70][131], Harray[71][131], Harray[72][131], Harray[73][131], Harray[74][131], Harray[75][131], Harray[76][131], Harray[77][131], Harray[78][131], Harray[79][131], Harray[80][131], Harray[81][131], Harray[82][131], Harray[83][131], Harray[84][131], Harray[85][131], Harray[86][131], Harray[87][131], Harray[88][131], Harray[89][131], Harray[90][131], Harray[91][131], Harray[92][131], Harray[93][131], Harray[94][131], Harray[95][131], Harray[96][131], Harray[97][131], Harray[98][131], Harray[99][131], Harray[100][131], Harray[101][131], Harray[102][131], Harray[103][131], Harray[104][131], Harray[105][131], Harray[106][131], Harray[107][131], Harray[108][131], Harray[109][131], Harray[110][131], Harray[111][131], Harray[112][131], Harray[113][131], Harray[114][131], Harray[115][131], Harray[116][131], Harray[117][131], Harray[118][131], Harray[119][131], Harray[120][131], Harray[121][131], Harray[122][131], Harray[123][131], Harray[124][131], Harray[125][131], Harray[126][131], Harray[127][131]};
assign h_col_132 = {Harray[0][132], Harray[1][132], Harray[2][132], Harray[3][132], Harray[4][132], Harray[5][132], Harray[6][132], Harray[7][132], Harray[8][132], Harray[9][132], Harray[10][132], Harray[11][132], Harray[12][132], Harray[13][132], Harray[14][132], Harray[15][132], Harray[16][132], Harray[17][132], Harray[18][132], Harray[19][132], Harray[20][132], Harray[21][132], Harray[22][132], Harray[23][132], Harray[24][132], Harray[25][132], Harray[26][132], Harray[27][132], Harray[28][132], Harray[29][132], Harray[30][132], Harray[31][132], Harray[32][132], Harray[33][132], Harray[34][132], Harray[35][132], Harray[36][132], Harray[37][132], Harray[38][132], Harray[39][132], Harray[40][132], Harray[41][132], Harray[42][132], Harray[43][132], Harray[44][132], Harray[45][132], Harray[46][132], Harray[47][132], Harray[48][132], Harray[49][132], Harray[50][132], Harray[51][132], Harray[52][132], Harray[53][132], Harray[54][132], Harray[55][132], Harray[56][132], Harray[57][132], Harray[58][132], Harray[59][132], Harray[60][132], Harray[61][132], Harray[62][132], Harray[63][132], Harray[64][132], Harray[65][132], Harray[66][132], Harray[67][132], Harray[68][132], Harray[69][132], Harray[70][132], Harray[71][132], Harray[72][132], Harray[73][132], Harray[74][132], Harray[75][132], Harray[76][132], Harray[77][132], Harray[78][132], Harray[79][132], Harray[80][132], Harray[81][132], Harray[82][132], Harray[83][132], Harray[84][132], Harray[85][132], Harray[86][132], Harray[87][132], Harray[88][132], Harray[89][132], Harray[90][132], Harray[91][132], Harray[92][132], Harray[93][132], Harray[94][132], Harray[95][132], Harray[96][132], Harray[97][132], Harray[98][132], Harray[99][132], Harray[100][132], Harray[101][132], Harray[102][132], Harray[103][132], Harray[104][132], Harray[105][132], Harray[106][132], Harray[107][132], Harray[108][132], Harray[109][132], Harray[110][132], Harray[111][132], Harray[112][132], Harray[113][132], Harray[114][132], Harray[115][132], Harray[116][132], Harray[117][132], Harray[118][132], Harray[119][132], Harray[120][132], Harray[121][132], Harray[122][132], Harray[123][132], Harray[124][132], Harray[125][132], Harray[126][132], Harray[127][132]};
assign h_col_133 = {Harray[0][133], Harray[1][133], Harray[2][133], Harray[3][133], Harray[4][133], Harray[5][133], Harray[6][133], Harray[7][133], Harray[8][133], Harray[9][133], Harray[10][133], Harray[11][133], Harray[12][133], Harray[13][133], Harray[14][133], Harray[15][133], Harray[16][133], Harray[17][133], Harray[18][133], Harray[19][133], Harray[20][133], Harray[21][133], Harray[22][133], Harray[23][133], Harray[24][133], Harray[25][133], Harray[26][133], Harray[27][133], Harray[28][133], Harray[29][133], Harray[30][133], Harray[31][133], Harray[32][133], Harray[33][133], Harray[34][133], Harray[35][133], Harray[36][133], Harray[37][133], Harray[38][133], Harray[39][133], Harray[40][133], Harray[41][133], Harray[42][133], Harray[43][133], Harray[44][133], Harray[45][133], Harray[46][133], Harray[47][133], Harray[48][133], Harray[49][133], Harray[50][133], Harray[51][133], Harray[52][133], Harray[53][133], Harray[54][133], Harray[55][133], Harray[56][133], Harray[57][133], Harray[58][133], Harray[59][133], Harray[60][133], Harray[61][133], Harray[62][133], Harray[63][133], Harray[64][133], Harray[65][133], Harray[66][133], Harray[67][133], Harray[68][133], Harray[69][133], Harray[70][133], Harray[71][133], Harray[72][133], Harray[73][133], Harray[74][133], Harray[75][133], Harray[76][133], Harray[77][133], Harray[78][133], Harray[79][133], Harray[80][133], Harray[81][133], Harray[82][133], Harray[83][133], Harray[84][133], Harray[85][133], Harray[86][133], Harray[87][133], Harray[88][133], Harray[89][133], Harray[90][133], Harray[91][133], Harray[92][133], Harray[93][133], Harray[94][133], Harray[95][133], Harray[96][133], Harray[97][133], Harray[98][133], Harray[99][133], Harray[100][133], Harray[101][133], Harray[102][133], Harray[103][133], Harray[104][133], Harray[105][133], Harray[106][133], Harray[107][133], Harray[108][133], Harray[109][133], Harray[110][133], Harray[111][133], Harray[112][133], Harray[113][133], Harray[114][133], Harray[115][133], Harray[116][133], Harray[117][133], Harray[118][133], Harray[119][133], Harray[120][133], Harray[121][133], Harray[122][133], Harray[123][133], Harray[124][133], Harray[125][133], Harray[126][133], Harray[127][133]};
assign h_col_134 = {Harray[0][134], Harray[1][134], Harray[2][134], Harray[3][134], Harray[4][134], Harray[5][134], Harray[6][134], Harray[7][134], Harray[8][134], Harray[9][134], Harray[10][134], Harray[11][134], Harray[12][134], Harray[13][134], Harray[14][134], Harray[15][134], Harray[16][134], Harray[17][134], Harray[18][134], Harray[19][134], Harray[20][134], Harray[21][134], Harray[22][134], Harray[23][134], Harray[24][134], Harray[25][134], Harray[26][134], Harray[27][134], Harray[28][134], Harray[29][134], Harray[30][134], Harray[31][134], Harray[32][134], Harray[33][134], Harray[34][134], Harray[35][134], Harray[36][134], Harray[37][134], Harray[38][134], Harray[39][134], Harray[40][134], Harray[41][134], Harray[42][134], Harray[43][134], Harray[44][134], Harray[45][134], Harray[46][134], Harray[47][134], Harray[48][134], Harray[49][134], Harray[50][134], Harray[51][134], Harray[52][134], Harray[53][134], Harray[54][134], Harray[55][134], Harray[56][134], Harray[57][134], Harray[58][134], Harray[59][134], Harray[60][134], Harray[61][134], Harray[62][134], Harray[63][134], Harray[64][134], Harray[65][134], Harray[66][134], Harray[67][134], Harray[68][134], Harray[69][134], Harray[70][134], Harray[71][134], Harray[72][134], Harray[73][134], Harray[74][134], Harray[75][134], Harray[76][134], Harray[77][134], Harray[78][134], Harray[79][134], Harray[80][134], Harray[81][134], Harray[82][134], Harray[83][134], Harray[84][134], Harray[85][134], Harray[86][134], Harray[87][134], Harray[88][134], Harray[89][134], Harray[90][134], Harray[91][134], Harray[92][134], Harray[93][134], Harray[94][134], Harray[95][134], Harray[96][134], Harray[97][134], Harray[98][134], Harray[99][134], Harray[100][134], Harray[101][134], Harray[102][134], Harray[103][134], Harray[104][134], Harray[105][134], Harray[106][134], Harray[107][134], Harray[108][134], Harray[109][134], Harray[110][134], Harray[111][134], Harray[112][134], Harray[113][134], Harray[114][134], Harray[115][134], Harray[116][134], Harray[117][134], Harray[118][134], Harray[119][134], Harray[120][134], Harray[121][134], Harray[122][134], Harray[123][134], Harray[124][134], Harray[125][134], Harray[126][134], Harray[127][134]};
assign h_col_135 = {Harray[0][135], Harray[1][135], Harray[2][135], Harray[3][135], Harray[4][135], Harray[5][135], Harray[6][135], Harray[7][135], Harray[8][135], Harray[9][135], Harray[10][135], Harray[11][135], Harray[12][135], Harray[13][135], Harray[14][135], Harray[15][135], Harray[16][135], Harray[17][135], Harray[18][135], Harray[19][135], Harray[20][135], Harray[21][135], Harray[22][135], Harray[23][135], Harray[24][135], Harray[25][135], Harray[26][135], Harray[27][135], Harray[28][135], Harray[29][135], Harray[30][135], Harray[31][135], Harray[32][135], Harray[33][135], Harray[34][135], Harray[35][135], Harray[36][135], Harray[37][135], Harray[38][135], Harray[39][135], Harray[40][135], Harray[41][135], Harray[42][135], Harray[43][135], Harray[44][135], Harray[45][135], Harray[46][135], Harray[47][135], Harray[48][135], Harray[49][135], Harray[50][135], Harray[51][135], Harray[52][135], Harray[53][135], Harray[54][135], Harray[55][135], Harray[56][135], Harray[57][135], Harray[58][135], Harray[59][135], Harray[60][135], Harray[61][135], Harray[62][135], Harray[63][135], Harray[64][135], Harray[65][135], Harray[66][135], Harray[67][135], Harray[68][135], Harray[69][135], Harray[70][135], Harray[71][135], Harray[72][135], Harray[73][135], Harray[74][135], Harray[75][135], Harray[76][135], Harray[77][135], Harray[78][135], Harray[79][135], Harray[80][135], Harray[81][135], Harray[82][135], Harray[83][135], Harray[84][135], Harray[85][135], Harray[86][135], Harray[87][135], Harray[88][135], Harray[89][135], Harray[90][135], Harray[91][135], Harray[92][135], Harray[93][135], Harray[94][135], Harray[95][135], Harray[96][135], Harray[97][135], Harray[98][135], Harray[99][135], Harray[100][135], Harray[101][135], Harray[102][135], Harray[103][135], Harray[104][135], Harray[105][135], Harray[106][135], Harray[107][135], Harray[108][135], Harray[109][135], Harray[110][135], Harray[111][135], Harray[112][135], Harray[113][135], Harray[114][135], Harray[115][135], Harray[116][135], Harray[117][135], Harray[118][135], Harray[119][135], Harray[120][135], Harray[121][135], Harray[122][135], Harray[123][135], Harray[124][135], Harray[125][135], Harray[126][135], Harray[127][135]};
assign h_col_136 = {Harray[0][136], Harray[1][136], Harray[2][136], Harray[3][136], Harray[4][136], Harray[5][136], Harray[6][136], Harray[7][136], Harray[8][136], Harray[9][136], Harray[10][136], Harray[11][136], Harray[12][136], Harray[13][136], Harray[14][136], Harray[15][136], Harray[16][136], Harray[17][136], Harray[18][136], Harray[19][136], Harray[20][136], Harray[21][136], Harray[22][136], Harray[23][136], Harray[24][136], Harray[25][136], Harray[26][136], Harray[27][136], Harray[28][136], Harray[29][136], Harray[30][136], Harray[31][136], Harray[32][136], Harray[33][136], Harray[34][136], Harray[35][136], Harray[36][136], Harray[37][136], Harray[38][136], Harray[39][136], Harray[40][136], Harray[41][136], Harray[42][136], Harray[43][136], Harray[44][136], Harray[45][136], Harray[46][136], Harray[47][136], Harray[48][136], Harray[49][136], Harray[50][136], Harray[51][136], Harray[52][136], Harray[53][136], Harray[54][136], Harray[55][136], Harray[56][136], Harray[57][136], Harray[58][136], Harray[59][136], Harray[60][136], Harray[61][136], Harray[62][136], Harray[63][136], Harray[64][136], Harray[65][136], Harray[66][136], Harray[67][136], Harray[68][136], Harray[69][136], Harray[70][136], Harray[71][136], Harray[72][136], Harray[73][136], Harray[74][136], Harray[75][136], Harray[76][136], Harray[77][136], Harray[78][136], Harray[79][136], Harray[80][136], Harray[81][136], Harray[82][136], Harray[83][136], Harray[84][136], Harray[85][136], Harray[86][136], Harray[87][136], Harray[88][136], Harray[89][136], Harray[90][136], Harray[91][136], Harray[92][136], Harray[93][136], Harray[94][136], Harray[95][136], Harray[96][136], Harray[97][136], Harray[98][136], Harray[99][136], Harray[100][136], Harray[101][136], Harray[102][136], Harray[103][136], Harray[104][136], Harray[105][136], Harray[106][136], Harray[107][136], Harray[108][136], Harray[109][136], Harray[110][136], Harray[111][136], Harray[112][136], Harray[113][136], Harray[114][136], Harray[115][136], Harray[116][136], Harray[117][136], Harray[118][136], Harray[119][136], Harray[120][136], Harray[121][136], Harray[122][136], Harray[123][136], Harray[124][136], Harray[125][136], Harray[126][136], Harray[127][136]};
assign h_col_137 = {Harray[0][137], Harray[1][137], Harray[2][137], Harray[3][137], Harray[4][137], Harray[5][137], Harray[6][137], Harray[7][137], Harray[8][137], Harray[9][137], Harray[10][137], Harray[11][137], Harray[12][137], Harray[13][137], Harray[14][137], Harray[15][137], Harray[16][137], Harray[17][137], Harray[18][137], Harray[19][137], Harray[20][137], Harray[21][137], Harray[22][137], Harray[23][137], Harray[24][137], Harray[25][137], Harray[26][137], Harray[27][137], Harray[28][137], Harray[29][137], Harray[30][137], Harray[31][137], Harray[32][137], Harray[33][137], Harray[34][137], Harray[35][137], Harray[36][137], Harray[37][137], Harray[38][137], Harray[39][137], Harray[40][137], Harray[41][137], Harray[42][137], Harray[43][137], Harray[44][137], Harray[45][137], Harray[46][137], Harray[47][137], Harray[48][137], Harray[49][137], Harray[50][137], Harray[51][137], Harray[52][137], Harray[53][137], Harray[54][137], Harray[55][137], Harray[56][137], Harray[57][137], Harray[58][137], Harray[59][137], Harray[60][137], Harray[61][137], Harray[62][137], Harray[63][137], Harray[64][137], Harray[65][137], Harray[66][137], Harray[67][137], Harray[68][137], Harray[69][137], Harray[70][137], Harray[71][137], Harray[72][137], Harray[73][137], Harray[74][137], Harray[75][137], Harray[76][137], Harray[77][137], Harray[78][137], Harray[79][137], Harray[80][137], Harray[81][137], Harray[82][137], Harray[83][137], Harray[84][137], Harray[85][137], Harray[86][137], Harray[87][137], Harray[88][137], Harray[89][137], Harray[90][137], Harray[91][137], Harray[92][137], Harray[93][137], Harray[94][137], Harray[95][137], Harray[96][137], Harray[97][137], Harray[98][137], Harray[99][137], Harray[100][137], Harray[101][137], Harray[102][137], Harray[103][137], Harray[104][137], Harray[105][137], Harray[106][137], Harray[107][137], Harray[108][137], Harray[109][137], Harray[110][137], Harray[111][137], Harray[112][137], Harray[113][137], Harray[114][137], Harray[115][137], Harray[116][137], Harray[117][137], Harray[118][137], Harray[119][137], Harray[120][137], Harray[121][137], Harray[122][137], Harray[123][137], Harray[124][137], Harray[125][137], Harray[126][137], Harray[127][137]};
assign h_col_138 = {Harray[0][138], Harray[1][138], Harray[2][138], Harray[3][138], Harray[4][138], Harray[5][138], Harray[6][138], Harray[7][138], Harray[8][138], Harray[9][138], Harray[10][138], Harray[11][138], Harray[12][138], Harray[13][138], Harray[14][138], Harray[15][138], Harray[16][138], Harray[17][138], Harray[18][138], Harray[19][138], Harray[20][138], Harray[21][138], Harray[22][138], Harray[23][138], Harray[24][138], Harray[25][138], Harray[26][138], Harray[27][138], Harray[28][138], Harray[29][138], Harray[30][138], Harray[31][138], Harray[32][138], Harray[33][138], Harray[34][138], Harray[35][138], Harray[36][138], Harray[37][138], Harray[38][138], Harray[39][138], Harray[40][138], Harray[41][138], Harray[42][138], Harray[43][138], Harray[44][138], Harray[45][138], Harray[46][138], Harray[47][138], Harray[48][138], Harray[49][138], Harray[50][138], Harray[51][138], Harray[52][138], Harray[53][138], Harray[54][138], Harray[55][138], Harray[56][138], Harray[57][138], Harray[58][138], Harray[59][138], Harray[60][138], Harray[61][138], Harray[62][138], Harray[63][138], Harray[64][138], Harray[65][138], Harray[66][138], Harray[67][138], Harray[68][138], Harray[69][138], Harray[70][138], Harray[71][138], Harray[72][138], Harray[73][138], Harray[74][138], Harray[75][138], Harray[76][138], Harray[77][138], Harray[78][138], Harray[79][138], Harray[80][138], Harray[81][138], Harray[82][138], Harray[83][138], Harray[84][138], Harray[85][138], Harray[86][138], Harray[87][138], Harray[88][138], Harray[89][138], Harray[90][138], Harray[91][138], Harray[92][138], Harray[93][138], Harray[94][138], Harray[95][138], Harray[96][138], Harray[97][138], Harray[98][138], Harray[99][138], Harray[100][138], Harray[101][138], Harray[102][138], Harray[103][138], Harray[104][138], Harray[105][138], Harray[106][138], Harray[107][138], Harray[108][138], Harray[109][138], Harray[110][138], Harray[111][138], Harray[112][138], Harray[113][138], Harray[114][138], Harray[115][138], Harray[116][138], Harray[117][138], Harray[118][138], Harray[119][138], Harray[120][138], Harray[121][138], Harray[122][138], Harray[123][138], Harray[124][138], Harray[125][138], Harray[126][138], Harray[127][138]};
assign h_col_139 = {Harray[0][139], Harray[1][139], Harray[2][139], Harray[3][139], Harray[4][139], Harray[5][139], Harray[6][139], Harray[7][139], Harray[8][139], Harray[9][139], Harray[10][139], Harray[11][139], Harray[12][139], Harray[13][139], Harray[14][139], Harray[15][139], Harray[16][139], Harray[17][139], Harray[18][139], Harray[19][139], Harray[20][139], Harray[21][139], Harray[22][139], Harray[23][139], Harray[24][139], Harray[25][139], Harray[26][139], Harray[27][139], Harray[28][139], Harray[29][139], Harray[30][139], Harray[31][139], Harray[32][139], Harray[33][139], Harray[34][139], Harray[35][139], Harray[36][139], Harray[37][139], Harray[38][139], Harray[39][139], Harray[40][139], Harray[41][139], Harray[42][139], Harray[43][139], Harray[44][139], Harray[45][139], Harray[46][139], Harray[47][139], Harray[48][139], Harray[49][139], Harray[50][139], Harray[51][139], Harray[52][139], Harray[53][139], Harray[54][139], Harray[55][139], Harray[56][139], Harray[57][139], Harray[58][139], Harray[59][139], Harray[60][139], Harray[61][139], Harray[62][139], Harray[63][139], Harray[64][139], Harray[65][139], Harray[66][139], Harray[67][139], Harray[68][139], Harray[69][139], Harray[70][139], Harray[71][139], Harray[72][139], Harray[73][139], Harray[74][139], Harray[75][139], Harray[76][139], Harray[77][139], Harray[78][139], Harray[79][139], Harray[80][139], Harray[81][139], Harray[82][139], Harray[83][139], Harray[84][139], Harray[85][139], Harray[86][139], Harray[87][139], Harray[88][139], Harray[89][139], Harray[90][139], Harray[91][139], Harray[92][139], Harray[93][139], Harray[94][139], Harray[95][139], Harray[96][139], Harray[97][139], Harray[98][139], Harray[99][139], Harray[100][139], Harray[101][139], Harray[102][139], Harray[103][139], Harray[104][139], Harray[105][139], Harray[106][139], Harray[107][139], Harray[108][139], Harray[109][139], Harray[110][139], Harray[111][139], Harray[112][139], Harray[113][139], Harray[114][139], Harray[115][139], Harray[116][139], Harray[117][139], Harray[118][139], Harray[119][139], Harray[120][139], Harray[121][139], Harray[122][139], Harray[123][139], Harray[124][139], Harray[125][139], Harray[126][139], Harray[127][139]};
assign h_col_140 = {Harray[0][140], Harray[1][140], Harray[2][140], Harray[3][140], Harray[4][140], Harray[5][140], Harray[6][140], Harray[7][140], Harray[8][140], Harray[9][140], Harray[10][140], Harray[11][140], Harray[12][140], Harray[13][140], Harray[14][140], Harray[15][140], Harray[16][140], Harray[17][140], Harray[18][140], Harray[19][140], Harray[20][140], Harray[21][140], Harray[22][140], Harray[23][140], Harray[24][140], Harray[25][140], Harray[26][140], Harray[27][140], Harray[28][140], Harray[29][140], Harray[30][140], Harray[31][140], Harray[32][140], Harray[33][140], Harray[34][140], Harray[35][140], Harray[36][140], Harray[37][140], Harray[38][140], Harray[39][140], Harray[40][140], Harray[41][140], Harray[42][140], Harray[43][140], Harray[44][140], Harray[45][140], Harray[46][140], Harray[47][140], Harray[48][140], Harray[49][140], Harray[50][140], Harray[51][140], Harray[52][140], Harray[53][140], Harray[54][140], Harray[55][140], Harray[56][140], Harray[57][140], Harray[58][140], Harray[59][140], Harray[60][140], Harray[61][140], Harray[62][140], Harray[63][140], Harray[64][140], Harray[65][140], Harray[66][140], Harray[67][140], Harray[68][140], Harray[69][140], Harray[70][140], Harray[71][140], Harray[72][140], Harray[73][140], Harray[74][140], Harray[75][140], Harray[76][140], Harray[77][140], Harray[78][140], Harray[79][140], Harray[80][140], Harray[81][140], Harray[82][140], Harray[83][140], Harray[84][140], Harray[85][140], Harray[86][140], Harray[87][140], Harray[88][140], Harray[89][140], Harray[90][140], Harray[91][140], Harray[92][140], Harray[93][140], Harray[94][140], Harray[95][140], Harray[96][140], Harray[97][140], Harray[98][140], Harray[99][140], Harray[100][140], Harray[101][140], Harray[102][140], Harray[103][140], Harray[104][140], Harray[105][140], Harray[106][140], Harray[107][140], Harray[108][140], Harray[109][140], Harray[110][140], Harray[111][140], Harray[112][140], Harray[113][140], Harray[114][140], Harray[115][140], Harray[116][140], Harray[117][140], Harray[118][140], Harray[119][140], Harray[120][140], Harray[121][140], Harray[122][140], Harray[123][140], Harray[124][140], Harray[125][140], Harray[126][140], Harray[127][140]};
assign h_col_141 = {Harray[0][141], Harray[1][141], Harray[2][141], Harray[3][141], Harray[4][141], Harray[5][141], Harray[6][141], Harray[7][141], Harray[8][141], Harray[9][141], Harray[10][141], Harray[11][141], Harray[12][141], Harray[13][141], Harray[14][141], Harray[15][141], Harray[16][141], Harray[17][141], Harray[18][141], Harray[19][141], Harray[20][141], Harray[21][141], Harray[22][141], Harray[23][141], Harray[24][141], Harray[25][141], Harray[26][141], Harray[27][141], Harray[28][141], Harray[29][141], Harray[30][141], Harray[31][141], Harray[32][141], Harray[33][141], Harray[34][141], Harray[35][141], Harray[36][141], Harray[37][141], Harray[38][141], Harray[39][141], Harray[40][141], Harray[41][141], Harray[42][141], Harray[43][141], Harray[44][141], Harray[45][141], Harray[46][141], Harray[47][141], Harray[48][141], Harray[49][141], Harray[50][141], Harray[51][141], Harray[52][141], Harray[53][141], Harray[54][141], Harray[55][141], Harray[56][141], Harray[57][141], Harray[58][141], Harray[59][141], Harray[60][141], Harray[61][141], Harray[62][141], Harray[63][141], Harray[64][141], Harray[65][141], Harray[66][141], Harray[67][141], Harray[68][141], Harray[69][141], Harray[70][141], Harray[71][141], Harray[72][141], Harray[73][141], Harray[74][141], Harray[75][141], Harray[76][141], Harray[77][141], Harray[78][141], Harray[79][141], Harray[80][141], Harray[81][141], Harray[82][141], Harray[83][141], Harray[84][141], Harray[85][141], Harray[86][141], Harray[87][141], Harray[88][141], Harray[89][141], Harray[90][141], Harray[91][141], Harray[92][141], Harray[93][141], Harray[94][141], Harray[95][141], Harray[96][141], Harray[97][141], Harray[98][141], Harray[99][141], Harray[100][141], Harray[101][141], Harray[102][141], Harray[103][141], Harray[104][141], Harray[105][141], Harray[106][141], Harray[107][141], Harray[108][141], Harray[109][141], Harray[110][141], Harray[111][141], Harray[112][141], Harray[113][141], Harray[114][141], Harray[115][141], Harray[116][141], Harray[117][141], Harray[118][141], Harray[119][141], Harray[120][141], Harray[121][141], Harray[122][141], Harray[123][141], Harray[124][141], Harray[125][141], Harray[126][141], Harray[127][141]};
assign h_col_142 = {Harray[0][142], Harray[1][142], Harray[2][142], Harray[3][142], Harray[4][142], Harray[5][142], Harray[6][142], Harray[7][142], Harray[8][142], Harray[9][142], Harray[10][142], Harray[11][142], Harray[12][142], Harray[13][142], Harray[14][142], Harray[15][142], Harray[16][142], Harray[17][142], Harray[18][142], Harray[19][142], Harray[20][142], Harray[21][142], Harray[22][142], Harray[23][142], Harray[24][142], Harray[25][142], Harray[26][142], Harray[27][142], Harray[28][142], Harray[29][142], Harray[30][142], Harray[31][142], Harray[32][142], Harray[33][142], Harray[34][142], Harray[35][142], Harray[36][142], Harray[37][142], Harray[38][142], Harray[39][142], Harray[40][142], Harray[41][142], Harray[42][142], Harray[43][142], Harray[44][142], Harray[45][142], Harray[46][142], Harray[47][142], Harray[48][142], Harray[49][142], Harray[50][142], Harray[51][142], Harray[52][142], Harray[53][142], Harray[54][142], Harray[55][142], Harray[56][142], Harray[57][142], Harray[58][142], Harray[59][142], Harray[60][142], Harray[61][142], Harray[62][142], Harray[63][142], Harray[64][142], Harray[65][142], Harray[66][142], Harray[67][142], Harray[68][142], Harray[69][142], Harray[70][142], Harray[71][142], Harray[72][142], Harray[73][142], Harray[74][142], Harray[75][142], Harray[76][142], Harray[77][142], Harray[78][142], Harray[79][142], Harray[80][142], Harray[81][142], Harray[82][142], Harray[83][142], Harray[84][142], Harray[85][142], Harray[86][142], Harray[87][142], Harray[88][142], Harray[89][142], Harray[90][142], Harray[91][142], Harray[92][142], Harray[93][142], Harray[94][142], Harray[95][142], Harray[96][142], Harray[97][142], Harray[98][142], Harray[99][142], Harray[100][142], Harray[101][142], Harray[102][142], Harray[103][142], Harray[104][142], Harray[105][142], Harray[106][142], Harray[107][142], Harray[108][142], Harray[109][142], Harray[110][142], Harray[111][142], Harray[112][142], Harray[113][142], Harray[114][142], Harray[115][142], Harray[116][142], Harray[117][142], Harray[118][142], Harray[119][142], Harray[120][142], Harray[121][142], Harray[122][142], Harray[123][142], Harray[124][142], Harray[125][142], Harray[126][142], Harray[127][142]};
assign h_col_143 = {Harray[0][143], Harray[1][143], Harray[2][143], Harray[3][143], Harray[4][143], Harray[5][143], Harray[6][143], Harray[7][143], Harray[8][143], Harray[9][143], Harray[10][143], Harray[11][143], Harray[12][143], Harray[13][143], Harray[14][143], Harray[15][143], Harray[16][143], Harray[17][143], Harray[18][143], Harray[19][143], Harray[20][143], Harray[21][143], Harray[22][143], Harray[23][143], Harray[24][143], Harray[25][143], Harray[26][143], Harray[27][143], Harray[28][143], Harray[29][143], Harray[30][143], Harray[31][143], Harray[32][143], Harray[33][143], Harray[34][143], Harray[35][143], Harray[36][143], Harray[37][143], Harray[38][143], Harray[39][143], Harray[40][143], Harray[41][143], Harray[42][143], Harray[43][143], Harray[44][143], Harray[45][143], Harray[46][143], Harray[47][143], Harray[48][143], Harray[49][143], Harray[50][143], Harray[51][143], Harray[52][143], Harray[53][143], Harray[54][143], Harray[55][143], Harray[56][143], Harray[57][143], Harray[58][143], Harray[59][143], Harray[60][143], Harray[61][143], Harray[62][143], Harray[63][143], Harray[64][143], Harray[65][143], Harray[66][143], Harray[67][143], Harray[68][143], Harray[69][143], Harray[70][143], Harray[71][143], Harray[72][143], Harray[73][143], Harray[74][143], Harray[75][143], Harray[76][143], Harray[77][143], Harray[78][143], Harray[79][143], Harray[80][143], Harray[81][143], Harray[82][143], Harray[83][143], Harray[84][143], Harray[85][143], Harray[86][143], Harray[87][143], Harray[88][143], Harray[89][143], Harray[90][143], Harray[91][143], Harray[92][143], Harray[93][143], Harray[94][143], Harray[95][143], Harray[96][143], Harray[97][143], Harray[98][143], Harray[99][143], Harray[100][143], Harray[101][143], Harray[102][143], Harray[103][143], Harray[104][143], Harray[105][143], Harray[106][143], Harray[107][143], Harray[108][143], Harray[109][143], Harray[110][143], Harray[111][143], Harray[112][143], Harray[113][143], Harray[114][143], Harray[115][143], Harray[116][143], Harray[117][143], Harray[118][143], Harray[119][143], Harray[120][143], Harray[121][143], Harray[122][143], Harray[123][143], Harray[124][143], Harray[125][143], Harray[126][143], Harray[127][143]};
assign h_col_144 = {Harray[0][144], Harray[1][144], Harray[2][144], Harray[3][144], Harray[4][144], Harray[5][144], Harray[6][144], Harray[7][144], Harray[8][144], Harray[9][144], Harray[10][144], Harray[11][144], Harray[12][144], Harray[13][144], Harray[14][144], Harray[15][144], Harray[16][144], Harray[17][144], Harray[18][144], Harray[19][144], Harray[20][144], Harray[21][144], Harray[22][144], Harray[23][144], Harray[24][144], Harray[25][144], Harray[26][144], Harray[27][144], Harray[28][144], Harray[29][144], Harray[30][144], Harray[31][144], Harray[32][144], Harray[33][144], Harray[34][144], Harray[35][144], Harray[36][144], Harray[37][144], Harray[38][144], Harray[39][144], Harray[40][144], Harray[41][144], Harray[42][144], Harray[43][144], Harray[44][144], Harray[45][144], Harray[46][144], Harray[47][144], Harray[48][144], Harray[49][144], Harray[50][144], Harray[51][144], Harray[52][144], Harray[53][144], Harray[54][144], Harray[55][144], Harray[56][144], Harray[57][144], Harray[58][144], Harray[59][144], Harray[60][144], Harray[61][144], Harray[62][144], Harray[63][144], Harray[64][144], Harray[65][144], Harray[66][144], Harray[67][144], Harray[68][144], Harray[69][144], Harray[70][144], Harray[71][144], Harray[72][144], Harray[73][144], Harray[74][144], Harray[75][144], Harray[76][144], Harray[77][144], Harray[78][144], Harray[79][144], Harray[80][144], Harray[81][144], Harray[82][144], Harray[83][144], Harray[84][144], Harray[85][144], Harray[86][144], Harray[87][144], Harray[88][144], Harray[89][144], Harray[90][144], Harray[91][144], Harray[92][144], Harray[93][144], Harray[94][144], Harray[95][144], Harray[96][144], Harray[97][144], Harray[98][144], Harray[99][144], Harray[100][144], Harray[101][144], Harray[102][144], Harray[103][144], Harray[104][144], Harray[105][144], Harray[106][144], Harray[107][144], Harray[108][144], Harray[109][144], Harray[110][144], Harray[111][144], Harray[112][144], Harray[113][144], Harray[114][144], Harray[115][144], Harray[116][144], Harray[117][144], Harray[118][144], Harray[119][144], Harray[120][144], Harray[121][144], Harray[122][144], Harray[123][144], Harray[124][144], Harray[125][144], Harray[126][144], Harray[127][144]};
assign h_col_145 = {Harray[0][145], Harray[1][145], Harray[2][145], Harray[3][145], Harray[4][145], Harray[5][145], Harray[6][145], Harray[7][145], Harray[8][145], Harray[9][145], Harray[10][145], Harray[11][145], Harray[12][145], Harray[13][145], Harray[14][145], Harray[15][145], Harray[16][145], Harray[17][145], Harray[18][145], Harray[19][145], Harray[20][145], Harray[21][145], Harray[22][145], Harray[23][145], Harray[24][145], Harray[25][145], Harray[26][145], Harray[27][145], Harray[28][145], Harray[29][145], Harray[30][145], Harray[31][145], Harray[32][145], Harray[33][145], Harray[34][145], Harray[35][145], Harray[36][145], Harray[37][145], Harray[38][145], Harray[39][145], Harray[40][145], Harray[41][145], Harray[42][145], Harray[43][145], Harray[44][145], Harray[45][145], Harray[46][145], Harray[47][145], Harray[48][145], Harray[49][145], Harray[50][145], Harray[51][145], Harray[52][145], Harray[53][145], Harray[54][145], Harray[55][145], Harray[56][145], Harray[57][145], Harray[58][145], Harray[59][145], Harray[60][145], Harray[61][145], Harray[62][145], Harray[63][145], Harray[64][145], Harray[65][145], Harray[66][145], Harray[67][145], Harray[68][145], Harray[69][145], Harray[70][145], Harray[71][145], Harray[72][145], Harray[73][145], Harray[74][145], Harray[75][145], Harray[76][145], Harray[77][145], Harray[78][145], Harray[79][145], Harray[80][145], Harray[81][145], Harray[82][145], Harray[83][145], Harray[84][145], Harray[85][145], Harray[86][145], Harray[87][145], Harray[88][145], Harray[89][145], Harray[90][145], Harray[91][145], Harray[92][145], Harray[93][145], Harray[94][145], Harray[95][145], Harray[96][145], Harray[97][145], Harray[98][145], Harray[99][145], Harray[100][145], Harray[101][145], Harray[102][145], Harray[103][145], Harray[104][145], Harray[105][145], Harray[106][145], Harray[107][145], Harray[108][145], Harray[109][145], Harray[110][145], Harray[111][145], Harray[112][145], Harray[113][145], Harray[114][145], Harray[115][145], Harray[116][145], Harray[117][145], Harray[118][145], Harray[119][145], Harray[120][145], Harray[121][145], Harray[122][145], Harray[123][145], Harray[124][145], Harray[125][145], Harray[126][145], Harray[127][145]};
assign h_col_146 = {Harray[0][146], Harray[1][146], Harray[2][146], Harray[3][146], Harray[4][146], Harray[5][146], Harray[6][146], Harray[7][146], Harray[8][146], Harray[9][146], Harray[10][146], Harray[11][146], Harray[12][146], Harray[13][146], Harray[14][146], Harray[15][146], Harray[16][146], Harray[17][146], Harray[18][146], Harray[19][146], Harray[20][146], Harray[21][146], Harray[22][146], Harray[23][146], Harray[24][146], Harray[25][146], Harray[26][146], Harray[27][146], Harray[28][146], Harray[29][146], Harray[30][146], Harray[31][146], Harray[32][146], Harray[33][146], Harray[34][146], Harray[35][146], Harray[36][146], Harray[37][146], Harray[38][146], Harray[39][146], Harray[40][146], Harray[41][146], Harray[42][146], Harray[43][146], Harray[44][146], Harray[45][146], Harray[46][146], Harray[47][146], Harray[48][146], Harray[49][146], Harray[50][146], Harray[51][146], Harray[52][146], Harray[53][146], Harray[54][146], Harray[55][146], Harray[56][146], Harray[57][146], Harray[58][146], Harray[59][146], Harray[60][146], Harray[61][146], Harray[62][146], Harray[63][146], Harray[64][146], Harray[65][146], Harray[66][146], Harray[67][146], Harray[68][146], Harray[69][146], Harray[70][146], Harray[71][146], Harray[72][146], Harray[73][146], Harray[74][146], Harray[75][146], Harray[76][146], Harray[77][146], Harray[78][146], Harray[79][146], Harray[80][146], Harray[81][146], Harray[82][146], Harray[83][146], Harray[84][146], Harray[85][146], Harray[86][146], Harray[87][146], Harray[88][146], Harray[89][146], Harray[90][146], Harray[91][146], Harray[92][146], Harray[93][146], Harray[94][146], Harray[95][146], Harray[96][146], Harray[97][146], Harray[98][146], Harray[99][146], Harray[100][146], Harray[101][146], Harray[102][146], Harray[103][146], Harray[104][146], Harray[105][146], Harray[106][146], Harray[107][146], Harray[108][146], Harray[109][146], Harray[110][146], Harray[111][146], Harray[112][146], Harray[113][146], Harray[114][146], Harray[115][146], Harray[116][146], Harray[117][146], Harray[118][146], Harray[119][146], Harray[120][146], Harray[121][146], Harray[122][146], Harray[123][146], Harray[124][146], Harray[125][146], Harray[126][146], Harray[127][146]};
assign h_col_147 = {Harray[0][147], Harray[1][147], Harray[2][147], Harray[3][147], Harray[4][147], Harray[5][147], Harray[6][147], Harray[7][147], Harray[8][147], Harray[9][147], Harray[10][147], Harray[11][147], Harray[12][147], Harray[13][147], Harray[14][147], Harray[15][147], Harray[16][147], Harray[17][147], Harray[18][147], Harray[19][147], Harray[20][147], Harray[21][147], Harray[22][147], Harray[23][147], Harray[24][147], Harray[25][147], Harray[26][147], Harray[27][147], Harray[28][147], Harray[29][147], Harray[30][147], Harray[31][147], Harray[32][147], Harray[33][147], Harray[34][147], Harray[35][147], Harray[36][147], Harray[37][147], Harray[38][147], Harray[39][147], Harray[40][147], Harray[41][147], Harray[42][147], Harray[43][147], Harray[44][147], Harray[45][147], Harray[46][147], Harray[47][147], Harray[48][147], Harray[49][147], Harray[50][147], Harray[51][147], Harray[52][147], Harray[53][147], Harray[54][147], Harray[55][147], Harray[56][147], Harray[57][147], Harray[58][147], Harray[59][147], Harray[60][147], Harray[61][147], Harray[62][147], Harray[63][147], Harray[64][147], Harray[65][147], Harray[66][147], Harray[67][147], Harray[68][147], Harray[69][147], Harray[70][147], Harray[71][147], Harray[72][147], Harray[73][147], Harray[74][147], Harray[75][147], Harray[76][147], Harray[77][147], Harray[78][147], Harray[79][147], Harray[80][147], Harray[81][147], Harray[82][147], Harray[83][147], Harray[84][147], Harray[85][147], Harray[86][147], Harray[87][147], Harray[88][147], Harray[89][147], Harray[90][147], Harray[91][147], Harray[92][147], Harray[93][147], Harray[94][147], Harray[95][147], Harray[96][147], Harray[97][147], Harray[98][147], Harray[99][147], Harray[100][147], Harray[101][147], Harray[102][147], Harray[103][147], Harray[104][147], Harray[105][147], Harray[106][147], Harray[107][147], Harray[108][147], Harray[109][147], Harray[110][147], Harray[111][147], Harray[112][147], Harray[113][147], Harray[114][147], Harray[115][147], Harray[116][147], Harray[117][147], Harray[118][147], Harray[119][147], Harray[120][147], Harray[121][147], Harray[122][147], Harray[123][147], Harray[124][147], Harray[125][147], Harray[126][147], Harray[127][147]};
assign h_col_148 = {Harray[0][148], Harray[1][148], Harray[2][148], Harray[3][148], Harray[4][148], Harray[5][148], Harray[6][148], Harray[7][148], Harray[8][148], Harray[9][148], Harray[10][148], Harray[11][148], Harray[12][148], Harray[13][148], Harray[14][148], Harray[15][148], Harray[16][148], Harray[17][148], Harray[18][148], Harray[19][148], Harray[20][148], Harray[21][148], Harray[22][148], Harray[23][148], Harray[24][148], Harray[25][148], Harray[26][148], Harray[27][148], Harray[28][148], Harray[29][148], Harray[30][148], Harray[31][148], Harray[32][148], Harray[33][148], Harray[34][148], Harray[35][148], Harray[36][148], Harray[37][148], Harray[38][148], Harray[39][148], Harray[40][148], Harray[41][148], Harray[42][148], Harray[43][148], Harray[44][148], Harray[45][148], Harray[46][148], Harray[47][148], Harray[48][148], Harray[49][148], Harray[50][148], Harray[51][148], Harray[52][148], Harray[53][148], Harray[54][148], Harray[55][148], Harray[56][148], Harray[57][148], Harray[58][148], Harray[59][148], Harray[60][148], Harray[61][148], Harray[62][148], Harray[63][148], Harray[64][148], Harray[65][148], Harray[66][148], Harray[67][148], Harray[68][148], Harray[69][148], Harray[70][148], Harray[71][148], Harray[72][148], Harray[73][148], Harray[74][148], Harray[75][148], Harray[76][148], Harray[77][148], Harray[78][148], Harray[79][148], Harray[80][148], Harray[81][148], Harray[82][148], Harray[83][148], Harray[84][148], Harray[85][148], Harray[86][148], Harray[87][148], Harray[88][148], Harray[89][148], Harray[90][148], Harray[91][148], Harray[92][148], Harray[93][148], Harray[94][148], Harray[95][148], Harray[96][148], Harray[97][148], Harray[98][148], Harray[99][148], Harray[100][148], Harray[101][148], Harray[102][148], Harray[103][148], Harray[104][148], Harray[105][148], Harray[106][148], Harray[107][148], Harray[108][148], Harray[109][148], Harray[110][148], Harray[111][148], Harray[112][148], Harray[113][148], Harray[114][148], Harray[115][148], Harray[116][148], Harray[117][148], Harray[118][148], Harray[119][148], Harray[120][148], Harray[121][148], Harray[122][148], Harray[123][148], Harray[124][148], Harray[125][148], Harray[126][148], Harray[127][148]};
assign h_col_149 = {Harray[0][149], Harray[1][149], Harray[2][149], Harray[3][149], Harray[4][149], Harray[5][149], Harray[6][149], Harray[7][149], Harray[8][149], Harray[9][149], Harray[10][149], Harray[11][149], Harray[12][149], Harray[13][149], Harray[14][149], Harray[15][149], Harray[16][149], Harray[17][149], Harray[18][149], Harray[19][149], Harray[20][149], Harray[21][149], Harray[22][149], Harray[23][149], Harray[24][149], Harray[25][149], Harray[26][149], Harray[27][149], Harray[28][149], Harray[29][149], Harray[30][149], Harray[31][149], Harray[32][149], Harray[33][149], Harray[34][149], Harray[35][149], Harray[36][149], Harray[37][149], Harray[38][149], Harray[39][149], Harray[40][149], Harray[41][149], Harray[42][149], Harray[43][149], Harray[44][149], Harray[45][149], Harray[46][149], Harray[47][149], Harray[48][149], Harray[49][149], Harray[50][149], Harray[51][149], Harray[52][149], Harray[53][149], Harray[54][149], Harray[55][149], Harray[56][149], Harray[57][149], Harray[58][149], Harray[59][149], Harray[60][149], Harray[61][149], Harray[62][149], Harray[63][149], Harray[64][149], Harray[65][149], Harray[66][149], Harray[67][149], Harray[68][149], Harray[69][149], Harray[70][149], Harray[71][149], Harray[72][149], Harray[73][149], Harray[74][149], Harray[75][149], Harray[76][149], Harray[77][149], Harray[78][149], Harray[79][149], Harray[80][149], Harray[81][149], Harray[82][149], Harray[83][149], Harray[84][149], Harray[85][149], Harray[86][149], Harray[87][149], Harray[88][149], Harray[89][149], Harray[90][149], Harray[91][149], Harray[92][149], Harray[93][149], Harray[94][149], Harray[95][149], Harray[96][149], Harray[97][149], Harray[98][149], Harray[99][149], Harray[100][149], Harray[101][149], Harray[102][149], Harray[103][149], Harray[104][149], Harray[105][149], Harray[106][149], Harray[107][149], Harray[108][149], Harray[109][149], Harray[110][149], Harray[111][149], Harray[112][149], Harray[113][149], Harray[114][149], Harray[115][149], Harray[116][149], Harray[117][149], Harray[118][149], Harray[119][149], Harray[120][149], Harray[121][149], Harray[122][149], Harray[123][149], Harray[124][149], Harray[125][149], Harray[126][149], Harray[127][149]};
assign h_col_150 = {Harray[0][150], Harray[1][150], Harray[2][150], Harray[3][150], Harray[4][150], Harray[5][150], Harray[6][150], Harray[7][150], Harray[8][150], Harray[9][150], Harray[10][150], Harray[11][150], Harray[12][150], Harray[13][150], Harray[14][150], Harray[15][150], Harray[16][150], Harray[17][150], Harray[18][150], Harray[19][150], Harray[20][150], Harray[21][150], Harray[22][150], Harray[23][150], Harray[24][150], Harray[25][150], Harray[26][150], Harray[27][150], Harray[28][150], Harray[29][150], Harray[30][150], Harray[31][150], Harray[32][150], Harray[33][150], Harray[34][150], Harray[35][150], Harray[36][150], Harray[37][150], Harray[38][150], Harray[39][150], Harray[40][150], Harray[41][150], Harray[42][150], Harray[43][150], Harray[44][150], Harray[45][150], Harray[46][150], Harray[47][150], Harray[48][150], Harray[49][150], Harray[50][150], Harray[51][150], Harray[52][150], Harray[53][150], Harray[54][150], Harray[55][150], Harray[56][150], Harray[57][150], Harray[58][150], Harray[59][150], Harray[60][150], Harray[61][150], Harray[62][150], Harray[63][150], Harray[64][150], Harray[65][150], Harray[66][150], Harray[67][150], Harray[68][150], Harray[69][150], Harray[70][150], Harray[71][150], Harray[72][150], Harray[73][150], Harray[74][150], Harray[75][150], Harray[76][150], Harray[77][150], Harray[78][150], Harray[79][150], Harray[80][150], Harray[81][150], Harray[82][150], Harray[83][150], Harray[84][150], Harray[85][150], Harray[86][150], Harray[87][150], Harray[88][150], Harray[89][150], Harray[90][150], Harray[91][150], Harray[92][150], Harray[93][150], Harray[94][150], Harray[95][150], Harray[96][150], Harray[97][150], Harray[98][150], Harray[99][150], Harray[100][150], Harray[101][150], Harray[102][150], Harray[103][150], Harray[104][150], Harray[105][150], Harray[106][150], Harray[107][150], Harray[108][150], Harray[109][150], Harray[110][150], Harray[111][150], Harray[112][150], Harray[113][150], Harray[114][150], Harray[115][150], Harray[116][150], Harray[117][150], Harray[118][150], Harray[119][150], Harray[120][150], Harray[121][150], Harray[122][150], Harray[123][150], Harray[124][150], Harray[125][150], Harray[126][150], Harray[127][150]};
assign h_col_151 = {Harray[0][151], Harray[1][151], Harray[2][151], Harray[3][151], Harray[4][151], Harray[5][151], Harray[6][151], Harray[7][151], Harray[8][151], Harray[9][151], Harray[10][151], Harray[11][151], Harray[12][151], Harray[13][151], Harray[14][151], Harray[15][151], Harray[16][151], Harray[17][151], Harray[18][151], Harray[19][151], Harray[20][151], Harray[21][151], Harray[22][151], Harray[23][151], Harray[24][151], Harray[25][151], Harray[26][151], Harray[27][151], Harray[28][151], Harray[29][151], Harray[30][151], Harray[31][151], Harray[32][151], Harray[33][151], Harray[34][151], Harray[35][151], Harray[36][151], Harray[37][151], Harray[38][151], Harray[39][151], Harray[40][151], Harray[41][151], Harray[42][151], Harray[43][151], Harray[44][151], Harray[45][151], Harray[46][151], Harray[47][151], Harray[48][151], Harray[49][151], Harray[50][151], Harray[51][151], Harray[52][151], Harray[53][151], Harray[54][151], Harray[55][151], Harray[56][151], Harray[57][151], Harray[58][151], Harray[59][151], Harray[60][151], Harray[61][151], Harray[62][151], Harray[63][151], Harray[64][151], Harray[65][151], Harray[66][151], Harray[67][151], Harray[68][151], Harray[69][151], Harray[70][151], Harray[71][151], Harray[72][151], Harray[73][151], Harray[74][151], Harray[75][151], Harray[76][151], Harray[77][151], Harray[78][151], Harray[79][151], Harray[80][151], Harray[81][151], Harray[82][151], Harray[83][151], Harray[84][151], Harray[85][151], Harray[86][151], Harray[87][151], Harray[88][151], Harray[89][151], Harray[90][151], Harray[91][151], Harray[92][151], Harray[93][151], Harray[94][151], Harray[95][151], Harray[96][151], Harray[97][151], Harray[98][151], Harray[99][151], Harray[100][151], Harray[101][151], Harray[102][151], Harray[103][151], Harray[104][151], Harray[105][151], Harray[106][151], Harray[107][151], Harray[108][151], Harray[109][151], Harray[110][151], Harray[111][151], Harray[112][151], Harray[113][151], Harray[114][151], Harray[115][151], Harray[116][151], Harray[117][151], Harray[118][151], Harray[119][151], Harray[120][151], Harray[121][151], Harray[122][151], Harray[123][151], Harray[124][151], Harray[125][151], Harray[126][151], Harray[127][151]};
assign h_col_152 = {Harray[0][152], Harray[1][152], Harray[2][152], Harray[3][152], Harray[4][152], Harray[5][152], Harray[6][152], Harray[7][152], Harray[8][152], Harray[9][152], Harray[10][152], Harray[11][152], Harray[12][152], Harray[13][152], Harray[14][152], Harray[15][152], Harray[16][152], Harray[17][152], Harray[18][152], Harray[19][152], Harray[20][152], Harray[21][152], Harray[22][152], Harray[23][152], Harray[24][152], Harray[25][152], Harray[26][152], Harray[27][152], Harray[28][152], Harray[29][152], Harray[30][152], Harray[31][152], Harray[32][152], Harray[33][152], Harray[34][152], Harray[35][152], Harray[36][152], Harray[37][152], Harray[38][152], Harray[39][152], Harray[40][152], Harray[41][152], Harray[42][152], Harray[43][152], Harray[44][152], Harray[45][152], Harray[46][152], Harray[47][152], Harray[48][152], Harray[49][152], Harray[50][152], Harray[51][152], Harray[52][152], Harray[53][152], Harray[54][152], Harray[55][152], Harray[56][152], Harray[57][152], Harray[58][152], Harray[59][152], Harray[60][152], Harray[61][152], Harray[62][152], Harray[63][152], Harray[64][152], Harray[65][152], Harray[66][152], Harray[67][152], Harray[68][152], Harray[69][152], Harray[70][152], Harray[71][152], Harray[72][152], Harray[73][152], Harray[74][152], Harray[75][152], Harray[76][152], Harray[77][152], Harray[78][152], Harray[79][152], Harray[80][152], Harray[81][152], Harray[82][152], Harray[83][152], Harray[84][152], Harray[85][152], Harray[86][152], Harray[87][152], Harray[88][152], Harray[89][152], Harray[90][152], Harray[91][152], Harray[92][152], Harray[93][152], Harray[94][152], Harray[95][152], Harray[96][152], Harray[97][152], Harray[98][152], Harray[99][152], Harray[100][152], Harray[101][152], Harray[102][152], Harray[103][152], Harray[104][152], Harray[105][152], Harray[106][152], Harray[107][152], Harray[108][152], Harray[109][152], Harray[110][152], Harray[111][152], Harray[112][152], Harray[113][152], Harray[114][152], Harray[115][152], Harray[116][152], Harray[117][152], Harray[118][152], Harray[119][152], Harray[120][152], Harray[121][152], Harray[122][152], Harray[123][152], Harray[124][152], Harray[125][152], Harray[126][152], Harray[127][152]};
assign h_col_153 = {Harray[0][153], Harray[1][153], Harray[2][153], Harray[3][153], Harray[4][153], Harray[5][153], Harray[6][153], Harray[7][153], Harray[8][153], Harray[9][153], Harray[10][153], Harray[11][153], Harray[12][153], Harray[13][153], Harray[14][153], Harray[15][153], Harray[16][153], Harray[17][153], Harray[18][153], Harray[19][153], Harray[20][153], Harray[21][153], Harray[22][153], Harray[23][153], Harray[24][153], Harray[25][153], Harray[26][153], Harray[27][153], Harray[28][153], Harray[29][153], Harray[30][153], Harray[31][153], Harray[32][153], Harray[33][153], Harray[34][153], Harray[35][153], Harray[36][153], Harray[37][153], Harray[38][153], Harray[39][153], Harray[40][153], Harray[41][153], Harray[42][153], Harray[43][153], Harray[44][153], Harray[45][153], Harray[46][153], Harray[47][153], Harray[48][153], Harray[49][153], Harray[50][153], Harray[51][153], Harray[52][153], Harray[53][153], Harray[54][153], Harray[55][153], Harray[56][153], Harray[57][153], Harray[58][153], Harray[59][153], Harray[60][153], Harray[61][153], Harray[62][153], Harray[63][153], Harray[64][153], Harray[65][153], Harray[66][153], Harray[67][153], Harray[68][153], Harray[69][153], Harray[70][153], Harray[71][153], Harray[72][153], Harray[73][153], Harray[74][153], Harray[75][153], Harray[76][153], Harray[77][153], Harray[78][153], Harray[79][153], Harray[80][153], Harray[81][153], Harray[82][153], Harray[83][153], Harray[84][153], Harray[85][153], Harray[86][153], Harray[87][153], Harray[88][153], Harray[89][153], Harray[90][153], Harray[91][153], Harray[92][153], Harray[93][153], Harray[94][153], Harray[95][153], Harray[96][153], Harray[97][153], Harray[98][153], Harray[99][153], Harray[100][153], Harray[101][153], Harray[102][153], Harray[103][153], Harray[104][153], Harray[105][153], Harray[106][153], Harray[107][153], Harray[108][153], Harray[109][153], Harray[110][153], Harray[111][153], Harray[112][153], Harray[113][153], Harray[114][153], Harray[115][153], Harray[116][153], Harray[117][153], Harray[118][153], Harray[119][153], Harray[120][153], Harray[121][153], Harray[122][153], Harray[123][153], Harray[124][153], Harray[125][153], Harray[126][153], Harray[127][153]};
assign h_col_154 = {Harray[0][154], Harray[1][154], Harray[2][154], Harray[3][154], Harray[4][154], Harray[5][154], Harray[6][154], Harray[7][154], Harray[8][154], Harray[9][154], Harray[10][154], Harray[11][154], Harray[12][154], Harray[13][154], Harray[14][154], Harray[15][154], Harray[16][154], Harray[17][154], Harray[18][154], Harray[19][154], Harray[20][154], Harray[21][154], Harray[22][154], Harray[23][154], Harray[24][154], Harray[25][154], Harray[26][154], Harray[27][154], Harray[28][154], Harray[29][154], Harray[30][154], Harray[31][154], Harray[32][154], Harray[33][154], Harray[34][154], Harray[35][154], Harray[36][154], Harray[37][154], Harray[38][154], Harray[39][154], Harray[40][154], Harray[41][154], Harray[42][154], Harray[43][154], Harray[44][154], Harray[45][154], Harray[46][154], Harray[47][154], Harray[48][154], Harray[49][154], Harray[50][154], Harray[51][154], Harray[52][154], Harray[53][154], Harray[54][154], Harray[55][154], Harray[56][154], Harray[57][154], Harray[58][154], Harray[59][154], Harray[60][154], Harray[61][154], Harray[62][154], Harray[63][154], Harray[64][154], Harray[65][154], Harray[66][154], Harray[67][154], Harray[68][154], Harray[69][154], Harray[70][154], Harray[71][154], Harray[72][154], Harray[73][154], Harray[74][154], Harray[75][154], Harray[76][154], Harray[77][154], Harray[78][154], Harray[79][154], Harray[80][154], Harray[81][154], Harray[82][154], Harray[83][154], Harray[84][154], Harray[85][154], Harray[86][154], Harray[87][154], Harray[88][154], Harray[89][154], Harray[90][154], Harray[91][154], Harray[92][154], Harray[93][154], Harray[94][154], Harray[95][154], Harray[96][154], Harray[97][154], Harray[98][154], Harray[99][154], Harray[100][154], Harray[101][154], Harray[102][154], Harray[103][154], Harray[104][154], Harray[105][154], Harray[106][154], Harray[107][154], Harray[108][154], Harray[109][154], Harray[110][154], Harray[111][154], Harray[112][154], Harray[113][154], Harray[114][154], Harray[115][154], Harray[116][154], Harray[117][154], Harray[118][154], Harray[119][154], Harray[120][154], Harray[121][154], Harray[122][154], Harray[123][154], Harray[124][154], Harray[125][154], Harray[126][154], Harray[127][154]};
assign h_col_155 = {Harray[0][155], Harray[1][155], Harray[2][155], Harray[3][155], Harray[4][155], Harray[5][155], Harray[6][155], Harray[7][155], Harray[8][155], Harray[9][155], Harray[10][155], Harray[11][155], Harray[12][155], Harray[13][155], Harray[14][155], Harray[15][155], Harray[16][155], Harray[17][155], Harray[18][155], Harray[19][155], Harray[20][155], Harray[21][155], Harray[22][155], Harray[23][155], Harray[24][155], Harray[25][155], Harray[26][155], Harray[27][155], Harray[28][155], Harray[29][155], Harray[30][155], Harray[31][155], Harray[32][155], Harray[33][155], Harray[34][155], Harray[35][155], Harray[36][155], Harray[37][155], Harray[38][155], Harray[39][155], Harray[40][155], Harray[41][155], Harray[42][155], Harray[43][155], Harray[44][155], Harray[45][155], Harray[46][155], Harray[47][155], Harray[48][155], Harray[49][155], Harray[50][155], Harray[51][155], Harray[52][155], Harray[53][155], Harray[54][155], Harray[55][155], Harray[56][155], Harray[57][155], Harray[58][155], Harray[59][155], Harray[60][155], Harray[61][155], Harray[62][155], Harray[63][155], Harray[64][155], Harray[65][155], Harray[66][155], Harray[67][155], Harray[68][155], Harray[69][155], Harray[70][155], Harray[71][155], Harray[72][155], Harray[73][155], Harray[74][155], Harray[75][155], Harray[76][155], Harray[77][155], Harray[78][155], Harray[79][155], Harray[80][155], Harray[81][155], Harray[82][155], Harray[83][155], Harray[84][155], Harray[85][155], Harray[86][155], Harray[87][155], Harray[88][155], Harray[89][155], Harray[90][155], Harray[91][155], Harray[92][155], Harray[93][155], Harray[94][155], Harray[95][155], Harray[96][155], Harray[97][155], Harray[98][155], Harray[99][155], Harray[100][155], Harray[101][155], Harray[102][155], Harray[103][155], Harray[104][155], Harray[105][155], Harray[106][155], Harray[107][155], Harray[108][155], Harray[109][155], Harray[110][155], Harray[111][155], Harray[112][155], Harray[113][155], Harray[114][155], Harray[115][155], Harray[116][155], Harray[117][155], Harray[118][155], Harray[119][155], Harray[120][155], Harray[121][155], Harray[122][155], Harray[123][155], Harray[124][155], Harray[125][155], Harray[126][155], Harray[127][155]};
assign h_col_156 = {Harray[0][156], Harray[1][156], Harray[2][156], Harray[3][156], Harray[4][156], Harray[5][156], Harray[6][156], Harray[7][156], Harray[8][156], Harray[9][156], Harray[10][156], Harray[11][156], Harray[12][156], Harray[13][156], Harray[14][156], Harray[15][156], Harray[16][156], Harray[17][156], Harray[18][156], Harray[19][156], Harray[20][156], Harray[21][156], Harray[22][156], Harray[23][156], Harray[24][156], Harray[25][156], Harray[26][156], Harray[27][156], Harray[28][156], Harray[29][156], Harray[30][156], Harray[31][156], Harray[32][156], Harray[33][156], Harray[34][156], Harray[35][156], Harray[36][156], Harray[37][156], Harray[38][156], Harray[39][156], Harray[40][156], Harray[41][156], Harray[42][156], Harray[43][156], Harray[44][156], Harray[45][156], Harray[46][156], Harray[47][156], Harray[48][156], Harray[49][156], Harray[50][156], Harray[51][156], Harray[52][156], Harray[53][156], Harray[54][156], Harray[55][156], Harray[56][156], Harray[57][156], Harray[58][156], Harray[59][156], Harray[60][156], Harray[61][156], Harray[62][156], Harray[63][156], Harray[64][156], Harray[65][156], Harray[66][156], Harray[67][156], Harray[68][156], Harray[69][156], Harray[70][156], Harray[71][156], Harray[72][156], Harray[73][156], Harray[74][156], Harray[75][156], Harray[76][156], Harray[77][156], Harray[78][156], Harray[79][156], Harray[80][156], Harray[81][156], Harray[82][156], Harray[83][156], Harray[84][156], Harray[85][156], Harray[86][156], Harray[87][156], Harray[88][156], Harray[89][156], Harray[90][156], Harray[91][156], Harray[92][156], Harray[93][156], Harray[94][156], Harray[95][156], Harray[96][156], Harray[97][156], Harray[98][156], Harray[99][156], Harray[100][156], Harray[101][156], Harray[102][156], Harray[103][156], Harray[104][156], Harray[105][156], Harray[106][156], Harray[107][156], Harray[108][156], Harray[109][156], Harray[110][156], Harray[111][156], Harray[112][156], Harray[113][156], Harray[114][156], Harray[115][156], Harray[116][156], Harray[117][156], Harray[118][156], Harray[119][156], Harray[120][156], Harray[121][156], Harray[122][156], Harray[123][156], Harray[124][156], Harray[125][156], Harray[126][156], Harray[127][156]};
assign h_col_157 = {Harray[0][157], Harray[1][157], Harray[2][157], Harray[3][157], Harray[4][157], Harray[5][157], Harray[6][157], Harray[7][157], Harray[8][157], Harray[9][157], Harray[10][157], Harray[11][157], Harray[12][157], Harray[13][157], Harray[14][157], Harray[15][157], Harray[16][157], Harray[17][157], Harray[18][157], Harray[19][157], Harray[20][157], Harray[21][157], Harray[22][157], Harray[23][157], Harray[24][157], Harray[25][157], Harray[26][157], Harray[27][157], Harray[28][157], Harray[29][157], Harray[30][157], Harray[31][157], Harray[32][157], Harray[33][157], Harray[34][157], Harray[35][157], Harray[36][157], Harray[37][157], Harray[38][157], Harray[39][157], Harray[40][157], Harray[41][157], Harray[42][157], Harray[43][157], Harray[44][157], Harray[45][157], Harray[46][157], Harray[47][157], Harray[48][157], Harray[49][157], Harray[50][157], Harray[51][157], Harray[52][157], Harray[53][157], Harray[54][157], Harray[55][157], Harray[56][157], Harray[57][157], Harray[58][157], Harray[59][157], Harray[60][157], Harray[61][157], Harray[62][157], Harray[63][157], Harray[64][157], Harray[65][157], Harray[66][157], Harray[67][157], Harray[68][157], Harray[69][157], Harray[70][157], Harray[71][157], Harray[72][157], Harray[73][157], Harray[74][157], Harray[75][157], Harray[76][157], Harray[77][157], Harray[78][157], Harray[79][157], Harray[80][157], Harray[81][157], Harray[82][157], Harray[83][157], Harray[84][157], Harray[85][157], Harray[86][157], Harray[87][157], Harray[88][157], Harray[89][157], Harray[90][157], Harray[91][157], Harray[92][157], Harray[93][157], Harray[94][157], Harray[95][157], Harray[96][157], Harray[97][157], Harray[98][157], Harray[99][157], Harray[100][157], Harray[101][157], Harray[102][157], Harray[103][157], Harray[104][157], Harray[105][157], Harray[106][157], Harray[107][157], Harray[108][157], Harray[109][157], Harray[110][157], Harray[111][157], Harray[112][157], Harray[113][157], Harray[114][157], Harray[115][157], Harray[116][157], Harray[117][157], Harray[118][157], Harray[119][157], Harray[120][157], Harray[121][157], Harray[122][157], Harray[123][157], Harray[124][157], Harray[125][157], Harray[126][157], Harray[127][157]};
assign h_col_158 = {Harray[0][158], Harray[1][158], Harray[2][158], Harray[3][158], Harray[4][158], Harray[5][158], Harray[6][158], Harray[7][158], Harray[8][158], Harray[9][158], Harray[10][158], Harray[11][158], Harray[12][158], Harray[13][158], Harray[14][158], Harray[15][158], Harray[16][158], Harray[17][158], Harray[18][158], Harray[19][158], Harray[20][158], Harray[21][158], Harray[22][158], Harray[23][158], Harray[24][158], Harray[25][158], Harray[26][158], Harray[27][158], Harray[28][158], Harray[29][158], Harray[30][158], Harray[31][158], Harray[32][158], Harray[33][158], Harray[34][158], Harray[35][158], Harray[36][158], Harray[37][158], Harray[38][158], Harray[39][158], Harray[40][158], Harray[41][158], Harray[42][158], Harray[43][158], Harray[44][158], Harray[45][158], Harray[46][158], Harray[47][158], Harray[48][158], Harray[49][158], Harray[50][158], Harray[51][158], Harray[52][158], Harray[53][158], Harray[54][158], Harray[55][158], Harray[56][158], Harray[57][158], Harray[58][158], Harray[59][158], Harray[60][158], Harray[61][158], Harray[62][158], Harray[63][158], Harray[64][158], Harray[65][158], Harray[66][158], Harray[67][158], Harray[68][158], Harray[69][158], Harray[70][158], Harray[71][158], Harray[72][158], Harray[73][158], Harray[74][158], Harray[75][158], Harray[76][158], Harray[77][158], Harray[78][158], Harray[79][158], Harray[80][158], Harray[81][158], Harray[82][158], Harray[83][158], Harray[84][158], Harray[85][158], Harray[86][158], Harray[87][158], Harray[88][158], Harray[89][158], Harray[90][158], Harray[91][158], Harray[92][158], Harray[93][158], Harray[94][158], Harray[95][158], Harray[96][158], Harray[97][158], Harray[98][158], Harray[99][158], Harray[100][158], Harray[101][158], Harray[102][158], Harray[103][158], Harray[104][158], Harray[105][158], Harray[106][158], Harray[107][158], Harray[108][158], Harray[109][158], Harray[110][158], Harray[111][158], Harray[112][158], Harray[113][158], Harray[114][158], Harray[115][158], Harray[116][158], Harray[117][158], Harray[118][158], Harray[119][158], Harray[120][158], Harray[121][158], Harray[122][158], Harray[123][158], Harray[124][158], Harray[125][158], Harray[126][158], Harray[127][158]};
assign h_col_159 = {Harray[0][159], Harray[1][159], Harray[2][159], Harray[3][159], Harray[4][159], Harray[5][159], Harray[6][159], Harray[7][159], Harray[8][159], Harray[9][159], Harray[10][159], Harray[11][159], Harray[12][159], Harray[13][159], Harray[14][159], Harray[15][159], Harray[16][159], Harray[17][159], Harray[18][159], Harray[19][159], Harray[20][159], Harray[21][159], Harray[22][159], Harray[23][159], Harray[24][159], Harray[25][159], Harray[26][159], Harray[27][159], Harray[28][159], Harray[29][159], Harray[30][159], Harray[31][159], Harray[32][159], Harray[33][159], Harray[34][159], Harray[35][159], Harray[36][159], Harray[37][159], Harray[38][159], Harray[39][159], Harray[40][159], Harray[41][159], Harray[42][159], Harray[43][159], Harray[44][159], Harray[45][159], Harray[46][159], Harray[47][159], Harray[48][159], Harray[49][159], Harray[50][159], Harray[51][159], Harray[52][159], Harray[53][159], Harray[54][159], Harray[55][159], Harray[56][159], Harray[57][159], Harray[58][159], Harray[59][159], Harray[60][159], Harray[61][159], Harray[62][159], Harray[63][159], Harray[64][159], Harray[65][159], Harray[66][159], Harray[67][159], Harray[68][159], Harray[69][159], Harray[70][159], Harray[71][159], Harray[72][159], Harray[73][159], Harray[74][159], Harray[75][159], Harray[76][159], Harray[77][159], Harray[78][159], Harray[79][159], Harray[80][159], Harray[81][159], Harray[82][159], Harray[83][159], Harray[84][159], Harray[85][159], Harray[86][159], Harray[87][159], Harray[88][159], Harray[89][159], Harray[90][159], Harray[91][159], Harray[92][159], Harray[93][159], Harray[94][159], Harray[95][159], Harray[96][159], Harray[97][159], Harray[98][159], Harray[99][159], Harray[100][159], Harray[101][159], Harray[102][159], Harray[103][159], Harray[104][159], Harray[105][159], Harray[106][159], Harray[107][159], Harray[108][159], Harray[109][159], Harray[110][159], Harray[111][159], Harray[112][159], Harray[113][159], Harray[114][159], Harray[115][159], Harray[116][159], Harray[117][159], Harray[118][159], Harray[119][159], Harray[120][159], Harray[121][159], Harray[122][159], Harray[123][159], Harray[124][159], Harray[125][159], Harray[126][159], Harray[127][159]};
assign h_col_160 = {Harray[0][160], Harray[1][160], Harray[2][160], Harray[3][160], Harray[4][160], Harray[5][160], Harray[6][160], Harray[7][160], Harray[8][160], Harray[9][160], Harray[10][160], Harray[11][160], Harray[12][160], Harray[13][160], Harray[14][160], Harray[15][160], Harray[16][160], Harray[17][160], Harray[18][160], Harray[19][160], Harray[20][160], Harray[21][160], Harray[22][160], Harray[23][160], Harray[24][160], Harray[25][160], Harray[26][160], Harray[27][160], Harray[28][160], Harray[29][160], Harray[30][160], Harray[31][160], Harray[32][160], Harray[33][160], Harray[34][160], Harray[35][160], Harray[36][160], Harray[37][160], Harray[38][160], Harray[39][160], Harray[40][160], Harray[41][160], Harray[42][160], Harray[43][160], Harray[44][160], Harray[45][160], Harray[46][160], Harray[47][160], Harray[48][160], Harray[49][160], Harray[50][160], Harray[51][160], Harray[52][160], Harray[53][160], Harray[54][160], Harray[55][160], Harray[56][160], Harray[57][160], Harray[58][160], Harray[59][160], Harray[60][160], Harray[61][160], Harray[62][160], Harray[63][160], Harray[64][160], Harray[65][160], Harray[66][160], Harray[67][160], Harray[68][160], Harray[69][160], Harray[70][160], Harray[71][160], Harray[72][160], Harray[73][160], Harray[74][160], Harray[75][160], Harray[76][160], Harray[77][160], Harray[78][160], Harray[79][160], Harray[80][160], Harray[81][160], Harray[82][160], Harray[83][160], Harray[84][160], Harray[85][160], Harray[86][160], Harray[87][160], Harray[88][160], Harray[89][160], Harray[90][160], Harray[91][160], Harray[92][160], Harray[93][160], Harray[94][160], Harray[95][160], Harray[96][160], Harray[97][160], Harray[98][160], Harray[99][160], Harray[100][160], Harray[101][160], Harray[102][160], Harray[103][160], Harray[104][160], Harray[105][160], Harray[106][160], Harray[107][160], Harray[108][160], Harray[109][160], Harray[110][160], Harray[111][160], Harray[112][160], Harray[113][160], Harray[114][160], Harray[115][160], Harray[116][160], Harray[117][160], Harray[118][160], Harray[119][160], Harray[120][160], Harray[121][160], Harray[122][160], Harray[123][160], Harray[124][160], Harray[125][160], Harray[126][160], Harray[127][160]};
assign h_col_161 = {Harray[0][161], Harray[1][161], Harray[2][161], Harray[3][161], Harray[4][161], Harray[5][161], Harray[6][161], Harray[7][161], Harray[8][161], Harray[9][161], Harray[10][161], Harray[11][161], Harray[12][161], Harray[13][161], Harray[14][161], Harray[15][161], Harray[16][161], Harray[17][161], Harray[18][161], Harray[19][161], Harray[20][161], Harray[21][161], Harray[22][161], Harray[23][161], Harray[24][161], Harray[25][161], Harray[26][161], Harray[27][161], Harray[28][161], Harray[29][161], Harray[30][161], Harray[31][161], Harray[32][161], Harray[33][161], Harray[34][161], Harray[35][161], Harray[36][161], Harray[37][161], Harray[38][161], Harray[39][161], Harray[40][161], Harray[41][161], Harray[42][161], Harray[43][161], Harray[44][161], Harray[45][161], Harray[46][161], Harray[47][161], Harray[48][161], Harray[49][161], Harray[50][161], Harray[51][161], Harray[52][161], Harray[53][161], Harray[54][161], Harray[55][161], Harray[56][161], Harray[57][161], Harray[58][161], Harray[59][161], Harray[60][161], Harray[61][161], Harray[62][161], Harray[63][161], Harray[64][161], Harray[65][161], Harray[66][161], Harray[67][161], Harray[68][161], Harray[69][161], Harray[70][161], Harray[71][161], Harray[72][161], Harray[73][161], Harray[74][161], Harray[75][161], Harray[76][161], Harray[77][161], Harray[78][161], Harray[79][161], Harray[80][161], Harray[81][161], Harray[82][161], Harray[83][161], Harray[84][161], Harray[85][161], Harray[86][161], Harray[87][161], Harray[88][161], Harray[89][161], Harray[90][161], Harray[91][161], Harray[92][161], Harray[93][161], Harray[94][161], Harray[95][161], Harray[96][161], Harray[97][161], Harray[98][161], Harray[99][161], Harray[100][161], Harray[101][161], Harray[102][161], Harray[103][161], Harray[104][161], Harray[105][161], Harray[106][161], Harray[107][161], Harray[108][161], Harray[109][161], Harray[110][161], Harray[111][161], Harray[112][161], Harray[113][161], Harray[114][161], Harray[115][161], Harray[116][161], Harray[117][161], Harray[118][161], Harray[119][161], Harray[120][161], Harray[121][161], Harray[122][161], Harray[123][161], Harray[124][161], Harray[125][161], Harray[126][161], Harray[127][161]};
assign h_col_162 = {Harray[0][162], Harray[1][162], Harray[2][162], Harray[3][162], Harray[4][162], Harray[5][162], Harray[6][162], Harray[7][162], Harray[8][162], Harray[9][162], Harray[10][162], Harray[11][162], Harray[12][162], Harray[13][162], Harray[14][162], Harray[15][162], Harray[16][162], Harray[17][162], Harray[18][162], Harray[19][162], Harray[20][162], Harray[21][162], Harray[22][162], Harray[23][162], Harray[24][162], Harray[25][162], Harray[26][162], Harray[27][162], Harray[28][162], Harray[29][162], Harray[30][162], Harray[31][162], Harray[32][162], Harray[33][162], Harray[34][162], Harray[35][162], Harray[36][162], Harray[37][162], Harray[38][162], Harray[39][162], Harray[40][162], Harray[41][162], Harray[42][162], Harray[43][162], Harray[44][162], Harray[45][162], Harray[46][162], Harray[47][162], Harray[48][162], Harray[49][162], Harray[50][162], Harray[51][162], Harray[52][162], Harray[53][162], Harray[54][162], Harray[55][162], Harray[56][162], Harray[57][162], Harray[58][162], Harray[59][162], Harray[60][162], Harray[61][162], Harray[62][162], Harray[63][162], Harray[64][162], Harray[65][162], Harray[66][162], Harray[67][162], Harray[68][162], Harray[69][162], Harray[70][162], Harray[71][162], Harray[72][162], Harray[73][162], Harray[74][162], Harray[75][162], Harray[76][162], Harray[77][162], Harray[78][162], Harray[79][162], Harray[80][162], Harray[81][162], Harray[82][162], Harray[83][162], Harray[84][162], Harray[85][162], Harray[86][162], Harray[87][162], Harray[88][162], Harray[89][162], Harray[90][162], Harray[91][162], Harray[92][162], Harray[93][162], Harray[94][162], Harray[95][162], Harray[96][162], Harray[97][162], Harray[98][162], Harray[99][162], Harray[100][162], Harray[101][162], Harray[102][162], Harray[103][162], Harray[104][162], Harray[105][162], Harray[106][162], Harray[107][162], Harray[108][162], Harray[109][162], Harray[110][162], Harray[111][162], Harray[112][162], Harray[113][162], Harray[114][162], Harray[115][162], Harray[116][162], Harray[117][162], Harray[118][162], Harray[119][162], Harray[120][162], Harray[121][162], Harray[122][162], Harray[123][162], Harray[124][162], Harray[125][162], Harray[126][162], Harray[127][162]};
assign h_col_163 = {Harray[0][163], Harray[1][163], Harray[2][163], Harray[3][163], Harray[4][163], Harray[5][163], Harray[6][163], Harray[7][163], Harray[8][163], Harray[9][163], Harray[10][163], Harray[11][163], Harray[12][163], Harray[13][163], Harray[14][163], Harray[15][163], Harray[16][163], Harray[17][163], Harray[18][163], Harray[19][163], Harray[20][163], Harray[21][163], Harray[22][163], Harray[23][163], Harray[24][163], Harray[25][163], Harray[26][163], Harray[27][163], Harray[28][163], Harray[29][163], Harray[30][163], Harray[31][163], Harray[32][163], Harray[33][163], Harray[34][163], Harray[35][163], Harray[36][163], Harray[37][163], Harray[38][163], Harray[39][163], Harray[40][163], Harray[41][163], Harray[42][163], Harray[43][163], Harray[44][163], Harray[45][163], Harray[46][163], Harray[47][163], Harray[48][163], Harray[49][163], Harray[50][163], Harray[51][163], Harray[52][163], Harray[53][163], Harray[54][163], Harray[55][163], Harray[56][163], Harray[57][163], Harray[58][163], Harray[59][163], Harray[60][163], Harray[61][163], Harray[62][163], Harray[63][163], Harray[64][163], Harray[65][163], Harray[66][163], Harray[67][163], Harray[68][163], Harray[69][163], Harray[70][163], Harray[71][163], Harray[72][163], Harray[73][163], Harray[74][163], Harray[75][163], Harray[76][163], Harray[77][163], Harray[78][163], Harray[79][163], Harray[80][163], Harray[81][163], Harray[82][163], Harray[83][163], Harray[84][163], Harray[85][163], Harray[86][163], Harray[87][163], Harray[88][163], Harray[89][163], Harray[90][163], Harray[91][163], Harray[92][163], Harray[93][163], Harray[94][163], Harray[95][163], Harray[96][163], Harray[97][163], Harray[98][163], Harray[99][163], Harray[100][163], Harray[101][163], Harray[102][163], Harray[103][163], Harray[104][163], Harray[105][163], Harray[106][163], Harray[107][163], Harray[108][163], Harray[109][163], Harray[110][163], Harray[111][163], Harray[112][163], Harray[113][163], Harray[114][163], Harray[115][163], Harray[116][163], Harray[117][163], Harray[118][163], Harray[119][163], Harray[120][163], Harray[121][163], Harray[122][163], Harray[123][163], Harray[124][163], Harray[125][163], Harray[126][163], Harray[127][163]};
assign h_col_164 = {Harray[0][164], Harray[1][164], Harray[2][164], Harray[3][164], Harray[4][164], Harray[5][164], Harray[6][164], Harray[7][164], Harray[8][164], Harray[9][164], Harray[10][164], Harray[11][164], Harray[12][164], Harray[13][164], Harray[14][164], Harray[15][164], Harray[16][164], Harray[17][164], Harray[18][164], Harray[19][164], Harray[20][164], Harray[21][164], Harray[22][164], Harray[23][164], Harray[24][164], Harray[25][164], Harray[26][164], Harray[27][164], Harray[28][164], Harray[29][164], Harray[30][164], Harray[31][164], Harray[32][164], Harray[33][164], Harray[34][164], Harray[35][164], Harray[36][164], Harray[37][164], Harray[38][164], Harray[39][164], Harray[40][164], Harray[41][164], Harray[42][164], Harray[43][164], Harray[44][164], Harray[45][164], Harray[46][164], Harray[47][164], Harray[48][164], Harray[49][164], Harray[50][164], Harray[51][164], Harray[52][164], Harray[53][164], Harray[54][164], Harray[55][164], Harray[56][164], Harray[57][164], Harray[58][164], Harray[59][164], Harray[60][164], Harray[61][164], Harray[62][164], Harray[63][164], Harray[64][164], Harray[65][164], Harray[66][164], Harray[67][164], Harray[68][164], Harray[69][164], Harray[70][164], Harray[71][164], Harray[72][164], Harray[73][164], Harray[74][164], Harray[75][164], Harray[76][164], Harray[77][164], Harray[78][164], Harray[79][164], Harray[80][164], Harray[81][164], Harray[82][164], Harray[83][164], Harray[84][164], Harray[85][164], Harray[86][164], Harray[87][164], Harray[88][164], Harray[89][164], Harray[90][164], Harray[91][164], Harray[92][164], Harray[93][164], Harray[94][164], Harray[95][164], Harray[96][164], Harray[97][164], Harray[98][164], Harray[99][164], Harray[100][164], Harray[101][164], Harray[102][164], Harray[103][164], Harray[104][164], Harray[105][164], Harray[106][164], Harray[107][164], Harray[108][164], Harray[109][164], Harray[110][164], Harray[111][164], Harray[112][164], Harray[113][164], Harray[114][164], Harray[115][164], Harray[116][164], Harray[117][164], Harray[118][164], Harray[119][164], Harray[120][164], Harray[121][164], Harray[122][164], Harray[123][164], Harray[124][164], Harray[125][164], Harray[126][164], Harray[127][164]};
assign h_col_165 = {Harray[0][165], Harray[1][165], Harray[2][165], Harray[3][165], Harray[4][165], Harray[5][165], Harray[6][165], Harray[7][165], Harray[8][165], Harray[9][165], Harray[10][165], Harray[11][165], Harray[12][165], Harray[13][165], Harray[14][165], Harray[15][165], Harray[16][165], Harray[17][165], Harray[18][165], Harray[19][165], Harray[20][165], Harray[21][165], Harray[22][165], Harray[23][165], Harray[24][165], Harray[25][165], Harray[26][165], Harray[27][165], Harray[28][165], Harray[29][165], Harray[30][165], Harray[31][165], Harray[32][165], Harray[33][165], Harray[34][165], Harray[35][165], Harray[36][165], Harray[37][165], Harray[38][165], Harray[39][165], Harray[40][165], Harray[41][165], Harray[42][165], Harray[43][165], Harray[44][165], Harray[45][165], Harray[46][165], Harray[47][165], Harray[48][165], Harray[49][165], Harray[50][165], Harray[51][165], Harray[52][165], Harray[53][165], Harray[54][165], Harray[55][165], Harray[56][165], Harray[57][165], Harray[58][165], Harray[59][165], Harray[60][165], Harray[61][165], Harray[62][165], Harray[63][165], Harray[64][165], Harray[65][165], Harray[66][165], Harray[67][165], Harray[68][165], Harray[69][165], Harray[70][165], Harray[71][165], Harray[72][165], Harray[73][165], Harray[74][165], Harray[75][165], Harray[76][165], Harray[77][165], Harray[78][165], Harray[79][165], Harray[80][165], Harray[81][165], Harray[82][165], Harray[83][165], Harray[84][165], Harray[85][165], Harray[86][165], Harray[87][165], Harray[88][165], Harray[89][165], Harray[90][165], Harray[91][165], Harray[92][165], Harray[93][165], Harray[94][165], Harray[95][165], Harray[96][165], Harray[97][165], Harray[98][165], Harray[99][165], Harray[100][165], Harray[101][165], Harray[102][165], Harray[103][165], Harray[104][165], Harray[105][165], Harray[106][165], Harray[107][165], Harray[108][165], Harray[109][165], Harray[110][165], Harray[111][165], Harray[112][165], Harray[113][165], Harray[114][165], Harray[115][165], Harray[116][165], Harray[117][165], Harray[118][165], Harray[119][165], Harray[120][165], Harray[121][165], Harray[122][165], Harray[123][165], Harray[124][165], Harray[125][165], Harray[126][165], Harray[127][165]};
assign h_col_166 = {Harray[0][166], Harray[1][166], Harray[2][166], Harray[3][166], Harray[4][166], Harray[5][166], Harray[6][166], Harray[7][166], Harray[8][166], Harray[9][166], Harray[10][166], Harray[11][166], Harray[12][166], Harray[13][166], Harray[14][166], Harray[15][166], Harray[16][166], Harray[17][166], Harray[18][166], Harray[19][166], Harray[20][166], Harray[21][166], Harray[22][166], Harray[23][166], Harray[24][166], Harray[25][166], Harray[26][166], Harray[27][166], Harray[28][166], Harray[29][166], Harray[30][166], Harray[31][166], Harray[32][166], Harray[33][166], Harray[34][166], Harray[35][166], Harray[36][166], Harray[37][166], Harray[38][166], Harray[39][166], Harray[40][166], Harray[41][166], Harray[42][166], Harray[43][166], Harray[44][166], Harray[45][166], Harray[46][166], Harray[47][166], Harray[48][166], Harray[49][166], Harray[50][166], Harray[51][166], Harray[52][166], Harray[53][166], Harray[54][166], Harray[55][166], Harray[56][166], Harray[57][166], Harray[58][166], Harray[59][166], Harray[60][166], Harray[61][166], Harray[62][166], Harray[63][166], Harray[64][166], Harray[65][166], Harray[66][166], Harray[67][166], Harray[68][166], Harray[69][166], Harray[70][166], Harray[71][166], Harray[72][166], Harray[73][166], Harray[74][166], Harray[75][166], Harray[76][166], Harray[77][166], Harray[78][166], Harray[79][166], Harray[80][166], Harray[81][166], Harray[82][166], Harray[83][166], Harray[84][166], Harray[85][166], Harray[86][166], Harray[87][166], Harray[88][166], Harray[89][166], Harray[90][166], Harray[91][166], Harray[92][166], Harray[93][166], Harray[94][166], Harray[95][166], Harray[96][166], Harray[97][166], Harray[98][166], Harray[99][166], Harray[100][166], Harray[101][166], Harray[102][166], Harray[103][166], Harray[104][166], Harray[105][166], Harray[106][166], Harray[107][166], Harray[108][166], Harray[109][166], Harray[110][166], Harray[111][166], Harray[112][166], Harray[113][166], Harray[114][166], Harray[115][166], Harray[116][166], Harray[117][166], Harray[118][166], Harray[119][166], Harray[120][166], Harray[121][166], Harray[122][166], Harray[123][166], Harray[124][166], Harray[125][166], Harray[126][166], Harray[127][166]};
assign h_col_167 = {Harray[0][167], Harray[1][167], Harray[2][167], Harray[3][167], Harray[4][167], Harray[5][167], Harray[6][167], Harray[7][167], Harray[8][167], Harray[9][167], Harray[10][167], Harray[11][167], Harray[12][167], Harray[13][167], Harray[14][167], Harray[15][167], Harray[16][167], Harray[17][167], Harray[18][167], Harray[19][167], Harray[20][167], Harray[21][167], Harray[22][167], Harray[23][167], Harray[24][167], Harray[25][167], Harray[26][167], Harray[27][167], Harray[28][167], Harray[29][167], Harray[30][167], Harray[31][167], Harray[32][167], Harray[33][167], Harray[34][167], Harray[35][167], Harray[36][167], Harray[37][167], Harray[38][167], Harray[39][167], Harray[40][167], Harray[41][167], Harray[42][167], Harray[43][167], Harray[44][167], Harray[45][167], Harray[46][167], Harray[47][167], Harray[48][167], Harray[49][167], Harray[50][167], Harray[51][167], Harray[52][167], Harray[53][167], Harray[54][167], Harray[55][167], Harray[56][167], Harray[57][167], Harray[58][167], Harray[59][167], Harray[60][167], Harray[61][167], Harray[62][167], Harray[63][167], Harray[64][167], Harray[65][167], Harray[66][167], Harray[67][167], Harray[68][167], Harray[69][167], Harray[70][167], Harray[71][167], Harray[72][167], Harray[73][167], Harray[74][167], Harray[75][167], Harray[76][167], Harray[77][167], Harray[78][167], Harray[79][167], Harray[80][167], Harray[81][167], Harray[82][167], Harray[83][167], Harray[84][167], Harray[85][167], Harray[86][167], Harray[87][167], Harray[88][167], Harray[89][167], Harray[90][167], Harray[91][167], Harray[92][167], Harray[93][167], Harray[94][167], Harray[95][167], Harray[96][167], Harray[97][167], Harray[98][167], Harray[99][167], Harray[100][167], Harray[101][167], Harray[102][167], Harray[103][167], Harray[104][167], Harray[105][167], Harray[106][167], Harray[107][167], Harray[108][167], Harray[109][167], Harray[110][167], Harray[111][167], Harray[112][167], Harray[113][167], Harray[114][167], Harray[115][167], Harray[116][167], Harray[117][167], Harray[118][167], Harray[119][167], Harray[120][167], Harray[121][167], Harray[122][167], Harray[123][167], Harray[124][167], Harray[125][167], Harray[126][167], Harray[127][167]};
assign h_col_168 = {Harray[0][168], Harray[1][168], Harray[2][168], Harray[3][168], Harray[4][168], Harray[5][168], Harray[6][168], Harray[7][168], Harray[8][168], Harray[9][168], Harray[10][168], Harray[11][168], Harray[12][168], Harray[13][168], Harray[14][168], Harray[15][168], Harray[16][168], Harray[17][168], Harray[18][168], Harray[19][168], Harray[20][168], Harray[21][168], Harray[22][168], Harray[23][168], Harray[24][168], Harray[25][168], Harray[26][168], Harray[27][168], Harray[28][168], Harray[29][168], Harray[30][168], Harray[31][168], Harray[32][168], Harray[33][168], Harray[34][168], Harray[35][168], Harray[36][168], Harray[37][168], Harray[38][168], Harray[39][168], Harray[40][168], Harray[41][168], Harray[42][168], Harray[43][168], Harray[44][168], Harray[45][168], Harray[46][168], Harray[47][168], Harray[48][168], Harray[49][168], Harray[50][168], Harray[51][168], Harray[52][168], Harray[53][168], Harray[54][168], Harray[55][168], Harray[56][168], Harray[57][168], Harray[58][168], Harray[59][168], Harray[60][168], Harray[61][168], Harray[62][168], Harray[63][168], Harray[64][168], Harray[65][168], Harray[66][168], Harray[67][168], Harray[68][168], Harray[69][168], Harray[70][168], Harray[71][168], Harray[72][168], Harray[73][168], Harray[74][168], Harray[75][168], Harray[76][168], Harray[77][168], Harray[78][168], Harray[79][168], Harray[80][168], Harray[81][168], Harray[82][168], Harray[83][168], Harray[84][168], Harray[85][168], Harray[86][168], Harray[87][168], Harray[88][168], Harray[89][168], Harray[90][168], Harray[91][168], Harray[92][168], Harray[93][168], Harray[94][168], Harray[95][168], Harray[96][168], Harray[97][168], Harray[98][168], Harray[99][168], Harray[100][168], Harray[101][168], Harray[102][168], Harray[103][168], Harray[104][168], Harray[105][168], Harray[106][168], Harray[107][168], Harray[108][168], Harray[109][168], Harray[110][168], Harray[111][168], Harray[112][168], Harray[113][168], Harray[114][168], Harray[115][168], Harray[116][168], Harray[117][168], Harray[118][168], Harray[119][168], Harray[120][168], Harray[121][168], Harray[122][168], Harray[123][168], Harray[124][168], Harray[125][168], Harray[126][168], Harray[127][168]};
assign h_col_169 = {Harray[0][169], Harray[1][169], Harray[2][169], Harray[3][169], Harray[4][169], Harray[5][169], Harray[6][169], Harray[7][169], Harray[8][169], Harray[9][169], Harray[10][169], Harray[11][169], Harray[12][169], Harray[13][169], Harray[14][169], Harray[15][169], Harray[16][169], Harray[17][169], Harray[18][169], Harray[19][169], Harray[20][169], Harray[21][169], Harray[22][169], Harray[23][169], Harray[24][169], Harray[25][169], Harray[26][169], Harray[27][169], Harray[28][169], Harray[29][169], Harray[30][169], Harray[31][169], Harray[32][169], Harray[33][169], Harray[34][169], Harray[35][169], Harray[36][169], Harray[37][169], Harray[38][169], Harray[39][169], Harray[40][169], Harray[41][169], Harray[42][169], Harray[43][169], Harray[44][169], Harray[45][169], Harray[46][169], Harray[47][169], Harray[48][169], Harray[49][169], Harray[50][169], Harray[51][169], Harray[52][169], Harray[53][169], Harray[54][169], Harray[55][169], Harray[56][169], Harray[57][169], Harray[58][169], Harray[59][169], Harray[60][169], Harray[61][169], Harray[62][169], Harray[63][169], Harray[64][169], Harray[65][169], Harray[66][169], Harray[67][169], Harray[68][169], Harray[69][169], Harray[70][169], Harray[71][169], Harray[72][169], Harray[73][169], Harray[74][169], Harray[75][169], Harray[76][169], Harray[77][169], Harray[78][169], Harray[79][169], Harray[80][169], Harray[81][169], Harray[82][169], Harray[83][169], Harray[84][169], Harray[85][169], Harray[86][169], Harray[87][169], Harray[88][169], Harray[89][169], Harray[90][169], Harray[91][169], Harray[92][169], Harray[93][169], Harray[94][169], Harray[95][169], Harray[96][169], Harray[97][169], Harray[98][169], Harray[99][169], Harray[100][169], Harray[101][169], Harray[102][169], Harray[103][169], Harray[104][169], Harray[105][169], Harray[106][169], Harray[107][169], Harray[108][169], Harray[109][169], Harray[110][169], Harray[111][169], Harray[112][169], Harray[113][169], Harray[114][169], Harray[115][169], Harray[116][169], Harray[117][169], Harray[118][169], Harray[119][169], Harray[120][169], Harray[121][169], Harray[122][169], Harray[123][169], Harray[124][169], Harray[125][169], Harray[126][169], Harray[127][169]};
assign h_col_170 = {Harray[0][170], Harray[1][170], Harray[2][170], Harray[3][170], Harray[4][170], Harray[5][170], Harray[6][170], Harray[7][170], Harray[8][170], Harray[9][170], Harray[10][170], Harray[11][170], Harray[12][170], Harray[13][170], Harray[14][170], Harray[15][170], Harray[16][170], Harray[17][170], Harray[18][170], Harray[19][170], Harray[20][170], Harray[21][170], Harray[22][170], Harray[23][170], Harray[24][170], Harray[25][170], Harray[26][170], Harray[27][170], Harray[28][170], Harray[29][170], Harray[30][170], Harray[31][170], Harray[32][170], Harray[33][170], Harray[34][170], Harray[35][170], Harray[36][170], Harray[37][170], Harray[38][170], Harray[39][170], Harray[40][170], Harray[41][170], Harray[42][170], Harray[43][170], Harray[44][170], Harray[45][170], Harray[46][170], Harray[47][170], Harray[48][170], Harray[49][170], Harray[50][170], Harray[51][170], Harray[52][170], Harray[53][170], Harray[54][170], Harray[55][170], Harray[56][170], Harray[57][170], Harray[58][170], Harray[59][170], Harray[60][170], Harray[61][170], Harray[62][170], Harray[63][170], Harray[64][170], Harray[65][170], Harray[66][170], Harray[67][170], Harray[68][170], Harray[69][170], Harray[70][170], Harray[71][170], Harray[72][170], Harray[73][170], Harray[74][170], Harray[75][170], Harray[76][170], Harray[77][170], Harray[78][170], Harray[79][170], Harray[80][170], Harray[81][170], Harray[82][170], Harray[83][170], Harray[84][170], Harray[85][170], Harray[86][170], Harray[87][170], Harray[88][170], Harray[89][170], Harray[90][170], Harray[91][170], Harray[92][170], Harray[93][170], Harray[94][170], Harray[95][170], Harray[96][170], Harray[97][170], Harray[98][170], Harray[99][170], Harray[100][170], Harray[101][170], Harray[102][170], Harray[103][170], Harray[104][170], Harray[105][170], Harray[106][170], Harray[107][170], Harray[108][170], Harray[109][170], Harray[110][170], Harray[111][170], Harray[112][170], Harray[113][170], Harray[114][170], Harray[115][170], Harray[116][170], Harray[117][170], Harray[118][170], Harray[119][170], Harray[120][170], Harray[121][170], Harray[122][170], Harray[123][170], Harray[124][170], Harray[125][170], Harray[126][170], Harray[127][170]};
assign h_col_171 = {Harray[0][171], Harray[1][171], Harray[2][171], Harray[3][171], Harray[4][171], Harray[5][171], Harray[6][171], Harray[7][171], Harray[8][171], Harray[9][171], Harray[10][171], Harray[11][171], Harray[12][171], Harray[13][171], Harray[14][171], Harray[15][171], Harray[16][171], Harray[17][171], Harray[18][171], Harray[19][171], Harray[20][171], Harray[21][171], Harray[22][171], Harray[23][171], Harray[24][171], Harray[25][171], Harray[26][171], Harray[27][171], Harray[28][171], Harray[29][171], Harray[30][171], Harray[31][171], Harray[32][171], Harray[33][171], Harray[34][171], Harray[35][171], Harray[36][171], Harray[37][171], Harray[38][171], Harray[39][171], Harray[40][171], Harray[41][171], Harray[42][171], Harray[43][171], Harray[44][171], Harray[45][171], Harray[46][171], Harray[47][171], Harray[48][171], Harray[49][171], Harray[50][171], Harray[51][171], Harray[52][171], Harray[53][171], Harray[54][171], Harray[55][171], Harray[56][171], Harray[57][171], Harray[58][171], Harray[59][171], Harray[60][171], Harray[61][171], Harray[62][171], Harray[63][171], Harray[64][171], Harray[65][171], Harray[66][171], Harray[67][171], Harray[68][171], Harray[69][171], Harray[70][171], Harray[71][171], Harray[72][171], Harray[73][171], Harray[74][171], Harray[75][171], Harray[76][171], Harray[77][171], Harray[78][171], Harray[79][171], Harray[80][171], Harray[81][171], Harray[82][171], Harray[83][171], Harray[84][171], Harray[85][171], Harray[86][171], Harray[87][171], Harray[88][171], Harray[89][171], Harray[90][171], Harray[91][171], Harray[92][171], Harray[93][171], Harray[94][171], Harray[95][171], Harray[96][171], Harray[97][171], Harray[98][171], Harray[99][171], Harray[100][171], Harray[101][171], Harray[102][171], Harray[103][171], Harray[104][171], Harray[105][171], Harray[106][171], Harray[107][171], Harray[108][171], Harray[109][171], Harray[110][171], Harray[111][171], Harray[112][171], Harray[113][171], Harray[114][171], Harray[115][171], Harray[116][171], Harray[117][171], Harray[118][171], Harray[119][171], Harray[120][171], Harray[121][171], Harray[122][171], Harray[123][171], Harray[124][171], Harray[125][171], Harray[126][171], Harray[127][171]};
assign h_col_172 = {Harray[0][172], Harray[1][172], Harray[2][172], Harray[3][172], Harray[4][172], Harray[5][172], Harray[6][172], Harray[7][172], Harray[8][172], Harray[9][172], Harray[10][172], Harray[11][172], Harray[12][172], Harray[13][172], Harray[14][172], Harray[15][172], Harray[16][172], Harray[17][172], Harray[18][172], Harray[19][172], Harray[20][172], Harray[21][172], Harray[22][172], Harray[23][172], Harray[24][172], Harray[25][172], Harray[26][172], Harray[27][172], Harray[28][172], Harray[29][172], Harray[30][172], Harray[31][172], Harray[32][172], Harray[33][172], Harray[34][172], Harray[35][172], Harray[36][172], Harray[37][172], Harray[38][172], Harray[39][172], Harray[40][172], Harray[41][172], Harray[42][172], Harray[43][172], Harray[44][172], Harray[45][172], Harray[46][172], Harray[47][172], Harray[48][172], Harray[49][172], Harray[50][172], Harray[51][172], Harray[52][172], Harray[53][172], Harray[54][172], Harray[55][172], Harray[56][172], Harray[57][172], Harray[58][172], Harray[59][172], Harray[60][172], Harray[61][172], Harray[62][172], Harray[63][172], Harray[64][172], Harray[65][172], Harray[66][172], Harray[67][172], Harray[68][172], Harray[69][172], Harray[70][172], Harray[71][172], Harray[72][172], Harray[73][172], Harray[74][172], Harray[75][172], Harray[76][172], Harray[77][172], Harray[78][172], Harray[79][172], Harray[80][172], Harray[81][172], Harray[82][172], Harray[83][172], Harray[84][172], Harray[85][172], Harray[86][172], Harray[87][172], Harray[88][172], Harray[89][172], Harray[90][172], Harray[91][172], Harray[92][172], Harray[93][172], Harray[94][172], Harray[95][172], Harray[96][172], Harray[97][172], Harray[98][172], Harray[99][172], Harray[100][172], Harray[101][172], Harray[102][172], Harray[103][172], Harray[104][172], Harray[105][172], Harray[106][172], Harray[107][172], Harray[108][172], Harray[109][172], Harray[110][172], Harray[111][172], Harray[112][172], Harray[113][172], Harray[114][172], Harray[115][172], Harray[116][172], Harray[117][172], Harray[118][172], Harray[119][172], Harray[120][172], Harray[121][172], Harray[122][172], Harray[123][172], Harray[124][172], Harray[125][172], Harray[126][172], Harray[127][172]};
assign h_col_173 = {Harray[0][173], Harray[1][173], Harray[2][173], Harray[3][173], Harray[4][173], Harray[5][173], Harray[6][173], Harray[7][173], Harray[8][173], Harray[9][173], Harray[10][173], Harray[11][173], Harray[12][173], Harray[13][173], Harray[14][173], Harray[15][173], Harray[16][173], Harray[17][173], Harray[18][173], Harray[19][173], Harray[20][173], Harray[21][173], Harray[22][173], Harray[23][173], Harray[24][173], Harray[25][173], Harray[26][173], Harray[27][173], Harray[28][173], Harray[29][173], Harray[30][173], Harray[31][173], Harray[32][173], Harray[33][173], Harray[34][173], Harray[35][173], Harray[36][173], Harray[37][173], Harray[38][173], Harray[39][173], Harray[40][173], Harray[41][173], Harray[42][173], Harray[43][173], Harray[44][173], Harray[45][173], Harray[46][173], Harray[47][173], Harray[48][173], Harray[49][173], Harray[50][173], Harray[51][173], Harray[52][173], Harray[53][173], Harray[54][173], Harray[55][173], Harray[56][173], Harray[57][173], Harray[58][173], Harray[59][173], Harray[60][173], Harray[61][173], Harray[62][173], Harray[63][173], Harray[64][173], Harray[65][173], Harray[66][173], Harray[67][173], Harray[68][173], Harray[69][173], Harray[70][173], Harray[71][173], Harray[72][173], Harray[73][173], Harray[74][173], Harray[75][173], Harray[76][173], Harray[77][173], Harray[78][173], Harray[79][173], Harray[80][173], Harray[81][173], Harray[82][173], Harray[83][173], Harray[84][173], Harray[85][173], Harray[86][173], Harray[87][173], Harray[88][173], Harray[89][173], Harray[90][173], Harray[91][173], Harray[92][173], Harray[93][173], Harray[94][173], Harray[95][173], Harray[96][173], Harray[97][173], Harray[98][173], Harray[99][173], Harray[100][173], Harray[101][173], Harray[102][173], Harray[103][173], Harray[104][173], Harray[105][173], Harray[106][173], Harray[107][173], Harray[108][173], Harray[109][173], Harray[110][173], Harray[111][173], Harray[112][173], Harray[113][173], Harray[114][173], Harray[115][173], Harray[116][173], Harray[117][173], Harray[118][173], Harray[119][173], Harray[120][173], Harray[121][173], Harray[122][173], Harray[123][173], Harray[124][173], Harray[125][173], Harray[126][173], Harray[127][173]};
assign h_col_174 = {Harray[0][174], Harray[1][174], Harray[2][174], Harray[3][174], Harray[4][174], Harray[5][174], Harray[6][174], Harray[7][174], Harray[8][174], Harray[9][174], Harray[10][174], Harray[11][174], Harray[12][174], Harray[13][174], Harray[14][174], Harray[15][174], Harray[16][174], Harray[17][174], Harray[18][174], Harray[19][174], Harray[20][174], Harray[21][174], Harray[22][174], Harray[23][174], Harray[24][174], Harray[25][174], Harray[26][174], Harray[27][174], Harray[28][174], Harray[29][174], Harray[30][174], Harray[31][174], Harray[32][174], Harray[33][174], Harray[34][174], Harray[35][174], Harray[36][174], Harray[37][174], Harray[38][174], Harray[39][174], Harray[40][174], Harray[41][174], Harray[42][174], Harray[43][174], Harray[44][174], Harray[45][174], Harray[46][174], Harray[47][174], Harray[48][174], Harray[49][174], Harray[50][174], Harray[51][174], Harray[52][174], Harray[53][174], Harray[54][174], Harray[55][174], Harray[56][174], Harray[57][174], Harray[58][174], Harray[59][174], Harray[60][174], Harray[61][174], Harray[62][174], Harray[63][174], Harray[64][174], Harray[65][174], Harray[66][174], Harray[67][174], Harray[68][174], Harray[69][174], Harray[70][174], Harray[71][174], Harray[72][174], Harray[73][174], Harray[74][174], Harray[75][174], Harray[76][174], Harray[77][174], Harray[78][174], Harray[79][174], Harray[80][174], Harray[81][174], Harray[82][174], Harray[83][174], Harray[84][174], Harray[85][174], Harray[86][174], Harray[87][174], Harray[88][174], Harray[89][174], Harray[90][174], Harray[91][174], Harray[92][174], Harray[93][174], Harray[94][174], Harray[95][174], Harray[96][174], Harray[97][174], Harray[98][174], Harray[99][174], Harray[100][174], Harray[101][174], Harray[102][174], Harray[103][174], Harray[104][174], Harray[105][174], Harray[106][174], Harray[107][174], Harray[108][174], Harray[109][174], Harray[110][174], Harray[111][174], Harray[112][174], Harray[113][174], Harray[114][174], Harray[115][174], Harray[116][174], Harray[117][174], Harray[118][174], Harray[119][174], Harray[120][174], Harray[121][174], Harray[122][174], Harray[123][174], Harray[124][174], Harray[125][174], Harray[126][174], Harray[127][174]};
assign h_col_175 = {Harray[0][175], Harray[1][175], Harray[2][175], Harray[3][175], Harray[4][175], Harray[5][175], Harray[6][175], Harray[7][175], Harray[8][175], Harray[9][175], Harray[10][175], Harray[11][175], Harray[12][175], Harray[13][175], Harray[14][175], Harray[15][175], Harray[16][175], Harray[17][175], Harray[18][175], Harray[19][175], Harray[20][175], Harray[21][175], Harray[22][175], Harray[23][175], Harray[24][175], Harray[25][175], Harray[26][175], Harray[27][175], Harray[28][175], Harray[29][175], Harray[30][175], Harray[31][175], Harray[32][175], Harray[33][175], Harray[34][175], Harray[35][175], Harray[36][175], Harray[37][175], Harray[38][175], Harray[39][175], Harray[40][175], Harray[41][175], Harray[42][175], Harray[43][175], Harray[44][175], Harray[45][175], Harray[46][175], Harray[47][175], Harray[48][175], Harray[49][175], Harray[50][175], Harray[51][175], Harray[52][175], Harray[53][175], Harray[54][175], Harray[55][175], Harray[56][175], Harray[57][175], Harray[58][175], Harray[59][175], Harray[60][175], Harray[61][175], Harray[62][175], Harray[63][175], Harray[64][175], Harray[65][175], Harray[66][175], Harray[67][175], Harray[68][175], Harray[69][175], Harray[70][175], Harray[71][175], Harray[72][175], Harray[73][175], Harray[74][175], Harray[75][175], Harray[76][175], Harray[77][175], Harray[78][175], Harray[79][175], Harray[80][175], Harray[81][175], Harray[82][175], Harray[83][175], Harray[84][175], Harray[85][175], Harray[86][175], Harray[87][175], Harray[88][175], Harray[89][175], Harray[90][175], Harray[91][175], Harray[92][175], Harray[93][175], Harray[94][175], Harray[95][175], Harray[96][175], Harray[97][175], Harray[98][175], Harray[99][175], Harray[100][175], Harray[101][175], Harray[102][175], Harray[103][175], Harray[104][175], Harray[105][175], Harray[106][175], Harray[107][175], Harray[108][175], Harray[109][175], Harray[110][175], Harray[111][175], Harray[112][175], Harray[113][175], Harray[114][175], Harray[115][175], Harray[116][175], Harray[117][175], Harray[118][175], Harray[119][175], Harray[120][175], Harray[121][175], Harray[122][175], Harray[123][175], Harray[124][175], Harray[125][175], Harray[126][175], Harray[127][175]};
assign h_col_176 = {Harray[0][176], Harray[1][176], Harray[2][176], Harray[3][176], Harray[4][176], Harray[5][176], Harray[6][176], Harray[7][176], Harray[8][176], Harray[9][176], Harray[10][176], Harray[11][176], Harray[12][176], Harray[13][176], Harray[14][176], Harray[15][176], Harray[16][176], Harray[17][176], Harray[18][176], Harray[19][176], Harray[20][176], Harray[21][176], Harray[22][176], Harray[23][176], Harray[24][176], Harray[25][176], Harray[26][176], Harray[27][176], Harray[28][176], Harray[29][176], Harray[30][176], Harray[31][176], Harray[32][176], Harray[33][176], Harray[34][176], Harray[35][176], Harray[36][176], Harray[37][176], Harray[38][176], Harray[39][176], Harray[40][176], Harray[41][176], Harray[42][176], Harray[43][176], Harray[44][176], Harray[45][176], Harray[46][176], Harray[47][176], Harray[48][176], Harray[49][176], Harray[50][176], Harray[51][176], Harray[52][176], Harray[53][176], Harray[54][176], Harray[55][176], Harray[56][176], Harray[57][176], Harray[58][176], Harray[59][176], Harray[60][176], Harray[61][176], Harray[62][176], Harray[63][176], Harray[64][176], Harray[65][176], Harray[66][176], Harray[67][176], Harray[68][176], Harray[69][176], Harray[70][176], Harray[71][176], Harray[72][176], Harray[73][176], Harray[74][176], Harray[75][176], Harray[76][176], Harray[77][176], Harray[78][176], Harray[79][176], Harray[80][176], Harray[81][176], Harray[82][176], Harray[83][176], Harray[84][176], Harray[85][176], Harray[86][176], Harray[87][176], Harray[88][176], Harray[89][176], Harray[90][176], Harray[91][176], Harray[92][176], Harray[93][176], Harray[94][176], Harray[95][176], Harray[96][176], Harray[97][176], Harray[98][176], Harray[99][176], Harray[100][176], Harray[101][176], Harray[102][176], Harray[103][176], Harray[104][176], Harray[105][176], Harray[106][176], Harray[107][176], Harray[108][176], Harray[109][176], Harray[110][176], Harray[111][176], Harray[112][176], Harray[113][176], Harray[114][176], Harray[115][176], Harray[116][176], Harray[117][176], Harray[118][176], Harray[119][176], Harray[120][176], Harray[121][176], Harray[122][176], Harray[123][176], Harray[124][176], Harray[125][176], Harray[126][176], Harray[127][176]};
assign h_col_177 = {Harray[0][177], Harray[1][177], Harray[2][177], Harray[3][177], Harray[4][177], Harray[5][177], Harray[6][177], Harray[7][177], Harray[8][177], Harray[9][177], Harray[10][177], Harray[11][177], Harray[12][177], Harray[13][177], Harray[14][177], Harray[15][177], Harray[16][177], Harray[17][177], Harray[18][177], Harray[19][177], Harray[20][177], Harray[21][177], Harray[22][177], Harray[23][177], Harray[24][177], Harray[25][177], Harray[26][177], Harray[27][177], Harray[28][177], Harray[29][177], Harray[30][177], Harray[31][177], Harray[32][177], Harray[33][177], Harray[34][177], Harray[35][177], Harray[36][177], Harray[37][177], Harray[38][177], Harray[39][177], Harray[40][177], Harray[41][177], Harray[42][177], Harray[43][177], Harray[44][177], Harray[45][177], Harray[46][177], Harray[47][177], Harray[48][177], Harray[49][177], Harray[50][177], Harray[51][177], Harray[52][177], Harray[53][177], Harray[54][177], Harray[55][177], Harray[56][177], Harray[57][177], Harray[58][177], Harray[59][177], Harray[60][177], Harray[61][177], Harray[62][177], Harray[63][177], Harray[64][177], Harray[65][177], Harray[66][177], Harray[67][177], Harray[68][177], Harray[69][177], Harray[70][177], Harray[71][177], Harray[72][177], Harray[73][177], Harray[74][177], Harray[75][177], Harray[76][177], Harray[77][177], Harray[78][177], Harray[79][177], Harray[80][177], Harray[81][177], Harray[82][177], Harray[83][177], Harray[84][177], Harray[85][177], Harray[86][177], Harray[87][177], Harray[88][177], Harray[89][177], Harray[90][177], Harray[91][177], Harray[92][177], Harray[93][177], Harray[94][177], Harray[95][177], Harray[96][177], Harray[97][177], Harray[98][177], Harray[99][177], Harray[100][177], Harray[101][177], Harray[102][177], Harray[103][177], Harray[104][177], Harray[105][177], Harray[106][177], Harray[107][177], Harray[108][177], Harray[109][177], Harray[110][177], Harray[111][177], Harray[112][177], Harray[113][177], Harray[114][177], Harray[115][177], Harray[116][177], Harray[117][177], Harray[118][177], Harray[119][177], Harray[120][177], Harray[121][177], Harray[122][177], Harray[123][177], Harray[124][177], Harray[125][177], Harray[126][177], Harray[127][177]};
assign h_col_178 = {Harray[0][178], Harray[1][178], Harray[2][178], Harray[3][178], Harray[4][178], Harray[5][178], Harray[6][178], Harray[7][178], Harray[8][178], Harray[9][178], Harray[10][178], Harray[11][178], Harray[12][178], Harray[13][178], Harray[14][178], Harray[15][178], Harray[16][178], Harray[17][178], Harray[18][178], Harray[19][178], Harray[20][178], Harray[21][178], Harray[22][178], Harray[23][178], Harray[24][178], Harray[25][178], Harray[26][178], Harray[27][178], Harray[28][178], Harray[29][178], Harray[30][178], Harray[31][178], Harray[32][178], Harray[33][178], Harray[34][178], Harray[35][178], Harray[36][178], Harray[37][178], Harray[38][178], Harray[39][178], Harray[40][178], Harray[41][178], Harray[42][178], Harray[43][178], Harray[44][178], Harray[45][178], Harray[46][178], Harray[47][178], Harray[48][178], Harray[49][178], Harray[50][178], Harray[51][178], Harray[52][178], Harray[53][178], Harray[54][178], Harray[55][178], Harray[56][178], Harray[57][178], Harray[58][178], Harray[59][178], Harray[60][178], Harray[61][178], Harray[62][178], Harray[63][178], Harray[64][178], Harray[65][178], Harray[66][178], Harray[67][178], Harray[68][178], Harray[69][178], Harray[70][178], Harray[71][178], Harray[72][178], Harray[73][178], Harray[74][178], Harray[75][178], Harray[76][178], Harray[77][178], Harray[78][178], Harray[79][178], Harray[80][178], Harray[81][178], Harray[82][178], Harray[83][178], Harray[84][178], Harray[85][178], Harray[86][178], Harray[87][178], Harray[88][178], Harray[89][178], Harray[90][178], Harray[91][178], Harray[92][178], Harray[93][178], Harray[94][178], Harray[95][178], Harray[96][178], Harray[97][178], Harray[98][178], Harray[99][178], Harray[100][178], Harray[101][178], Harray[102][178], Harray[103][178], Harray[104][178], Harray[105][178], Harray[106][178], Harray[107][178], Harray[108][178], Harray[109][178], Harray[110][178], Harray[111][178], Harray[112][178], Harray[113][178], Harray[114][178], Harray[115][178], Harray[116][178], Harray[117][178], Harray[118][178], Harray[119][178], Harray[120][178], Harray[121][178], Harray[122][178], Harray[123][178], Harray[124][178], Harray[125][178], Harray[126][178], Harray[127][178]};
assign h_col_179 = {Harray[0][179], Harray[1][179], Harray[2][179], Harray[3][179], Harray[4][179], Harray[5][179], Harray[6][179], Harray[7][179], Harray[8][179], Harray[9][179], Harray[10][179], Harray[11][179], Harray[12][179], Harray[13][179], Harray[14][179], Harray[15][179], Harray[16][179], Harray[17][179], Harray[18][179], Harray[19][179], Harray[20][179], Harray[21][179], Harray[22][179], Harray[23][179], Harray[24][179], Harray[25][179], Harray[26][179], Harray[27][179], Harray[28][179], Harray[29][179], Harray[30][179], Harray[31][179], Harray[32][179], Harray[33][179], Harray[34][179], Harray[35][179], Harray[36][179], Harray[37][179], Harray[38][179], Harray[39][179], Harray[40][179], Harray[41][179], Harray[42][179], Harray[43][179], Harray[44][179], Harray[45][179], Harray[46][179], Harray[47][179], Harray[48][179], Harray[49][179], Harray[50][179], Harray[51][179], Harray[52][179], Harray[53][179], Harray[54][179], Harray[55][179], Harray[56][179], Harray[57][179], Harray[58][179], Harray[59][179], Harray[60][179], Harray[61][179], Harray[62][179], Harray[63][179], Harray[64][179], Harray[65][179], Harray[66][179], Harray[67][179], Harray[68][179], Harray[69][179], Harray[70][179], Harray[71][179], Harray[72][179], Harray[73][179], Harray[74][179], Harray[75][179], Harray[76][179], Harray[77][179], Harray[78][179], Harray[79][179], Harray[80][179], Harray[81][179], Harray[82][179], Harray[83][179], Harray[84][179], Harray[85][179], Harray[86][179], Harray[87][179], Harray[88][179], Harray[89][179], Harray[90][179], Harray[91][179], Harray[92][179], Harray[93][179], Harray[94][179], Harray[95][179], Harray[96][179], Harray[97][179], Harray[98][179], Harray[99][179], Harray[100][179], Harray[101][179], Harray[102][179], Harray[103][179], Harray[104][179], Harray[105][179], Harray[106][179], Harray[107][179], Harray[108][179], Harray[109][179], Harray[110][179], Harray[111][179], Harray[112][179], Harray[113][179], Harray[114][179], Harray[115][179], Harray[116][179], Harray[117][179], Harray[118][179], Harray[119][179], Harray[120][179], Harray[121][179], Harray[122][179], Harray[123][179], Harray[124][179], Harray[125][179], Harray[126][179], Harray[127][179]};
assign h_col_180 = {Harray[0][180], Harray[1][180], Harray[2][180], Harray[3][180], Harray[4][180], Harray[5][180], Harray[6][180], Harray[7][180], Harray[8][180], Harray[9][180], Harray[10][180], Harray[11][180], Harray[12][180], Harray[13][180], Harray[14][180], Harray[15][180], Harray[16][180], Harray[17][180], Harray[18][180], Harray[19][180], Harray[20][180], Harray[21][180], Harray[22][180], Harray[23][180], Harray[24][180], Harray[25][180], Harray[26][180], Harray[27][180], Harray[28][180], Harray[29][180], Harray[30][180], Harray[31][180], Harray[32][180], Harray[33][180], Harray[34][180], Harray[35][180], Harray[36][180], Harray[37][180], Harray[38][180], Harray[39][180], Harray[40][180], Harray[41][180], Harray[42][180], Harray[43][180], Harray[44][180], Harray[45][180], Harray[46][180], Harray[47][180], Harray[48][180], Harray[49][180], Harray[50][180], Harray[51][180], Harray[52][180], Harray[53][180], Harray[54][180], Harray[55][180], Harray[56][180], Harray[57][180], Harray[58][180], Harray[59][180], Harray[60][180], Harray[61][180], Harray[62][180], Harray[63][180], Harray[64][180], Harray[65][180], Harray[66][180], Harray[67][180], Harray[68][180], Harray[69][180], Harray[70][180], Harray[71][180], Harray[72][180], Harray[73][180], Harray[74][180], Harray[75][180], Harray[76][180], Harray[77][180], Harray[78][180], Harray[79][180], Harray[80][180], Harray[81][180], Harray[82][180], Harray[83][180], Harray[84][180], Harray[85][180], Harray[86][180], Harray[87][180], Harray[88][180], Harray[89][180], Harray[90][180], Harray[91][180], Harray[92][180], Harray[93][180], Harray[94][180], Harray[95][180], Harray[96][180], Harray[97][180], Harray[98][180], Harray[99][180], Harray[100][180], Harray[101][180], Harray[102][180], Harray[103][180], Harray[104][180], Harray[105][180], Harray[106][180], Harray[107][180], Harray[108][180], Harray[109][180], Harray[110][180], Harray[111][180], Harray[112][180], Harray[113][180], Harray[114][180], Harray[115][180], Harray[116][180], Harray[117][180], Harray[118][180], Harray[119][180], Harray[120][180], Harray[121][180], Harray[122][180], Harray[123][180], Harray[124][180], Harray[125][180], Harray[126][180], Harray[127][180]};
assign h_col_181 = {Harray[0][181], Harray[1][181], Harray[2][181], Harray[3][181], Harray[4][181], Harray[5][181], Harray[6][181], Harray[7][181], Harray[8][181], Harray[9][181], Harray[10][181], Harray[11][181], Harray[12][181], Harray[13][181], Harray[14][181], Harray[15][181], Harray[16][181], Harray[17][181], Harray[18][181], Harray[19][181], Harray[20][181], Harray[21][181], Harray[22][181], Harray[23][181], Harray[24][181], Harray[25][181], Harray[26][181], Harray[27][181], Harray[28][181], Harray[29][181], Harray[30][181], Harray[31][181], Harray[32][181], Harray[33][181], Harray[34][181], Harray[35][181], Harray[36][181], Harray[37][181], Harray[38][181], Harray[39][181], Harray[40][181], Harray[41][181], Harray[42][181], Harray[43][181], Harray[44][181], Harray[45][181], Harray[46][181], Harray[47][181], Harray[48][181], Harray[49][181], Harray[50][181], Harray[51][181], Harray[52][181], Harray[53][181], Harray[54][181], Harray[55][181], Harray[56][181], Harray[57][181], Harray[58][181], Harray[59][181], Harray[60][181], Harray[61][181], Harray[62][181], Harray[63][181], Harray[64][181], Harray[65][181], Harray[66][181], Harray[67][181], Harray[68][181], Harray[69][181], Harray[70][181], Harray[71][181], Harray[72][181], Harray[73][181], Harray[74][181], Harray[75][181], Harray[76][181], Harray[77][181], Harray[78][181], Harray[79][181], Harray[80][181], Harray[81][181], Harray[82][181], Harray[83][181], Harray[84][181], Harray[85][181], Harray[86][181], Harray[87][181], Harray[88][181], Harray[89][181], Harray[90][181], Harray[91][181], Harray[92][181], Harray[93][181], Harray[94][181], Harray[95][181], Harray[96][181], Harray[97][181], Harray[98][181], Harray[99][181], Harray[100][181], Harray[101][181], Harray[102][181], Harray[103][181], Harray[104][181], Harray[105][181], Harray[106][181], Harray[107][181], Harray[108][181], Harray[109][181], Harray[110][181], Harray[111][181], Harray[112][181], Harray[113][181], Harray[114][181], Harray[115][181], Harray[116][181], Harray[117][181], Harray[118][181], Harray[119][181], Harray[120][181], Harray[121][181], Harray[122][181], Harray[123][181], Harray[124][181], Harray[125][181], Harray[126][181], Harray[127][181]};
assign h_col_182 = {Harray[0][182], Harray[1][182], Harray[2][182], Harray[3][182], Harray[4][182], Harray[5][182], Harray[6][182], Harray[7][182], Harray[8][182], Harray[9][182], Harray[10][182], Harray[11][182], Harray[12][182], Harray[13][182], Harray[14][182], Harray[15][182], Harray[16][182], Harray[17][182], Harray[18][182], Harray[19][182], Harray[20][182], Harray[21][182], Harray[22][182], Harray[23][182], Harray[24][182], Harray[25][182], Harray[26][182], Harray[27][182], Harray[28][182], Harray[29][182], Harray[30][182], Harray[31][182], Harray[32][182], Harray[33][182], Harray[34][182], Harray[35][182], Harray[36][182], Harray[37][182], Harray[38][182], Harray[39][182], Harray[40][182], Harray[41][182], Harray[42][182], Harray[43][182], Harray[44][182], Harray[45][182], Harray[46][182], Harray[47][182], Harray[48][182], Harray[49][182], Harray[50][182], Harray[51][182], Harray[52][182], Harray[53][182], Harray[54][182], Harray[55][182], Harray[56][182], Harray[57][182], Harray[58][182], Harray[59][182], Harray[60][182], Harray[61][182], Harray[62][182], Harray[63][182], Harray[64][182], Harray[65][182], Harray[66][182], Harray[67][182], Harray[68][182], Harray[69][182], Harray[70][182], Harray[71][182], Harray[72][182], Harray[73][182], Harray[74][182], Harray[75][182], Harray[76][182], Harray[77][182], Harray[78][182], Harray[79][182], Harray[80][182], Harray[81][182], Harray[82][182], Harray[83][182], Harray[84][182], Harray[85][182], Harray[86][182], Harray[87][182], Harray[88][182], Harray[89][182], Harray[90][182], Harray[91][182], Harray[92][182], Harray[93][182], Harray[94][182], Harray[95][182], Harray[96][182], Harray[97][182], Harray[98][182], Harray[99][182], Harray[100][182], Harray[101][182], Harray[102][182], Harray[103][182], Harray[104][182], Harray[105][182], Harray[106][182], Harray[107][182], Harray[108][182], Harray[109][182], Harray[110][182], Harray[111][182], Harray[112][182], Harray[113][182], Harray[114][182], Harray[115][182], Harray[116][182], Harray[117][182], Harray[118][182], Harray[119][182], Harray[120][182], Harray[121][182], Harray[122][182], Harray[123][182], Harray[124][182], Harray[125][182], Harray[126][182], Harray[127][182]};
assign h_col_183 = {Harray[0][183], Harray[1][183], Harray[2][183], Harray[3][183], Harray[4][183], Harray[5][183], Harray[6][183], Harray[7][183], Harray[8][183], Harray[9][183], Harray[10][183], Harray[11][183], Harray[12][183], Harray[13][183], Harray[14][183], Harray[15][183], Harray[16][183], Harray[17][183], Harray[18][183], Harray[19][183], Harray[20][183], Harray[21][183], Harray[22][183], Harray[23][183], Harray[24][183], Harray[25][183], Harray[26][183], Harray[27][183], Harray[28][183], Harray[29][183], Harray[30][183], Harray[31][183], Harray[32][183], Harray[33][183], Harray[34][183], Harray[35][183], Harray[36][183], Harray[37][183], Harray[38][183], Harray[39][183], Harray[40][183], Harray[41][183], Harray[42][183], Harray[43][183], Harray[44][183], Harray[45][183], Harray[46][183], Harray[47][183], Harray[48][183], Harray[49][183], Harray[50][183], Harray[51][183], Harray[52][183], Harray[53][183], Harray[54][183], Harray[55][183], Harray[56][183], Harray[57][183], Harray[58][183], Harray[59][183], Harray[60][183], Harray[61][183], Harray[62][183], Harray[63][183], Harray[64][183], Harray[65][183], Harray[66][183], Harray[67][183], Harray[68][183], Harray[69][183], Harray[70][183], Harray[71][183], Harray[72][183], Harray[73][183], Harray[74][183], Harray[75][183], Harray[76][183], Harray[77][183], Harray[78][183], Harray[79][183], Harray[80][183], Harray[81][183], Harray[82][183], Harray[83][183], Harray[84][183], Harray[85][183], Harray[86][183], Harray[87][183], Harray[88][183], Harray[89][183], Harray[90][183], Harray[91][183], Harray[92][183], Harray[93][183], Harray[94][183], Harray[95][183], Harray[96][183], Harray[97][183], Harray[98][183], Harray[99][183], Harray[100][183], Harray[101][183], Harray[102][183], Harray[103][183], Harray[104][183], Harray[105][183], Harray[106][183], Harray[107][183], Harray[108][183], Harray[109][183], Harray[110][183], Harray[111][183], Harray[112][183], Harray[113][183], Harray[114][183], Harray[115][183], Harray[116][183], Harray[117][183], Harray[118][183], Harray[119][183], Harray[120][183], Harray[121][183], Harray[122][183], Harray[123][183], Harray[124][183], Harray[125][183], Harray[126][183], Harray[127][183]};
assign h_col_184 = {Harray[0][184], Harray[1][184], Harray[2][184], Harray[3][184], Harray[4][184], Harray[5][184], Harray[6][184], Harray[7][184], Harray[8][184], Harray[9][184], Harray[10][184], Harray[11][184], Harray[12][184], Harray[13][184], Harray[14][184], Harray[15][184], Harray[16][184], Harray[17][184], Harray[18][184], Harray[19][184], Harray[20][184], Harray[21][184], Harray[22][184], Harray[23][184], Harray[24][184], Harray[25][184], Harray[26][184], Harray[27][184], Harray[28][184], Harray[29][184], Harray[30][184], Harray[31][184], Harray[32][184], Harray[33][184], Harray[34][184], Harray[35][184], Harray[36][184], Harray[37][184], Harray[38][184], Harray[39][184], Harray[40][184], Harray[41][184], Harray[42][184], Harray[43][184], Harray[44][184], Harray[45][184], Harray[46][184], Harray[47][184], Harray[48][184], Harray[49][184], Harray[50][184], Harray[51][184], Harray[52][184], Harray[53][184], Harray[54][184], Harray[55][184], Harray[56][184], Harray[57][184], Harray[58][184], Harray[59][184], Harray[60][184], Harray[61][184], Harray[62][184], Harray[63][184], Harray[64][184], Harray[65][184], Harray[66][184], Harray[67][184], Harray[68][184], Harray[69][184], Harray[70][184], Harray[71][184], Harray[72][184], Harray[73][184], Harray[74][184], Harray[75][184], Harray[76][184], Harray[77][184], Harray[78][184], Harray[79][184], Harray[80][184], Harray[81][184], Harray[82][184], Harray[83][184], Harray[84][184], Harray[85][184], Harray[86][184], Harray[87][184], Harray[88][184], Harray[89][184], Harray[90][184], Harray[91][184], Harray[92][184], Harray[93][184], Harray[94][184], Harray[95][184], Harray[96][184], Harray[97][184], Harray[98][184], Harray[99][184], Harray[100][184], Harray[101][184], Harray[102][184], Harray[103][184], Harray[104][184], Harray[105][184], Harray[106][184], Harray[107][184], Harray[108][184], Harray[109][184], Harray[110][184], Harray[111][184], Harray[112][184], Harray[113][184], Harray[114][184], Harray[115][184], Harray[116][184], Harray[117][184], Harray[118][184], Harray[119][184], Harray[120][184], Harray[121][184], Harray[122][184], Harray[123][184], Harray[124][184], Harray[125][184], Harray[126][184], Harray[127][184]};
assign h_col_185 = {Harray[0][185], Harray[1][185], Harray[2][185], Harray[3][185], Harray[4][185], Harray[5][185], Harray[6][185], Harray[7][185], Harray[8][185], Harray[9][185], Harray[10][185], Harray[11][185], Harray[12][185], Harray[13][185], Harray[14][185], Harray[15][185], Harray[16][185], Harray[17][185], Harray[18][185], Harray[19][185], Harray[20][185], Harray[21][185], Harray[22][185], Harray[23][185], Harray[24][185], Harray[25][185], Harray[26][185], Harray[27][185], Harray[28][185], Harray[29][185], Harray[30][185], Harray[31][185], Harray[32][185], Harray[33][185], Harray[34][185], Harray[35][185], Harray[36][185], Harray[37][185], Harray[38][185], Harray[39][185], Harray[40][185], Harray[41][185], Harray[42][185], Harray[43][185], Harray[44][185], Harray[45][185], Harray[46][185], Harray[47][185], Harray[48][185], Harray[49][185], Harray[50][185], Harray[51][185], Harray[52][185], Harray[53][185], Harray[54][185], Harray[55][185], Harray[56][185], Harray[57][185], Harray[58][185], Harray[59][185], Harray[60][185], Harray[61][185], Harray[62][185], Harray[63][185], Harray[64][185], Harray[65][185], Harray[66][185], Harray[67][185], Harray[68][185], Harray[69][185], Harray[70][185], Harray[71][185], Harray[72][185], Harray[73][185], Harray[74][185], Harray[75][185], Harray[76][185], Harray[77][185], Harray[78][185], Harray[79][185], Harray[80][185], Harray[81][185], Harray[82][185], Harray[83][185], Harray[84][185], Harray[85][185], Harray[86][185], Harray[87][185], Harray[88][185], Harray[89][185], Harray[90][185], Harray[91][185], Harray[92][185], Harray[93][185], Harray[94][185], Harray[95][185], Harray[96][185], Harray[97][185], Harray[98][185], Harray[99][185], Harray[100][185], Harray[101][185], Harray[102][185], Harray[103][185], Harray[104][185], Harray[105][185], Harray[106][185], Harray[107][185], Harray[108][185], Harray[109][185], Harray[110][185], Harray[111][185], Harray[112][185], Harray[113][185], Harray[114][185], Harray[115][185], Harray[116][185], Harray[117][185], Harray[118][185], Harray[119][185], Harray[120][185], Harray[121][185], Harray[122][185], Harray[123][185], Harray[124][185], Harray[125][185], Harray[126][185], Harray[127][185]};
assign h_col_186 = {Harray[0][186], Harray[1][186], Harray[2][186], Harray[3][186], Harray[4][186], Harray[5][186], Harray[6][186], Harray[7][186], Harray[8][186], Harray[9][186], Harray[10][186], Harray[11][186], Harray[12][186], Harray[13][186], Harray[14][186], Harray[15][186], Harray[16][186], Harray[17][186], Harray[18][186], Harray[19][186], Harray[20][186], Harray[21][186], Harray[22][186], Harray[23][186], Harray[24][186], Harray[25][186], Harray[26][186], Harray[27][186], Harray[28][186], Harray[29][186], Harray[30][186], Harray[31][186], Harray[32][186], Harray[33][186], Harray[34][186], Harray[35][186], Harray[36][186], Harray[37][186], Harray[38][186], Harray[39][186], Harray[40][186], Harray[41][186], Harray[42][186], Harray[43][186], Harray[44][186], Harray[45][186], Harray[46][186], Harray[47][186], Harray[48][186], Harray[49][186], Harray[50][186], Harray[51][186], Harray[52][186], Harray[53][186], Harray[54][186], Harray[55][186], Harray[56][186], Harray[57][186], Harray[58][186], Harray[59][186], Harray[60][186], Harray[61][186], Harray[62][186], Harray[63][186], Harray[64][186], Harray[65][186], Harray[66][186], Harray[67][186], Harray[68][186], Harray[69][186], Harray[70][186], Harray[71][186], Harray[72][186], Harray[73][186], Harray[74][186], Harray[75][186], Harray[76][186], Harray[77][186], Harray[78][186], Harray[79][186], Harray[80][186], Harray[81][186], Harray[82][186], Harray[83][186], Harray[84][186], Harray[85][186], Harray[86][186], Harray[87][186], Harray[88][186], Harray[89][186], Harray[90][186], Harray[91][186], Harray[92][186], Harray[93][186], Harray[94][186], Harray[95][186], Harray[96][186], Harray[97][186], Harray[98][186], Harray[99][186], Harray[100][186], Harray[101][186], Harray[102][186], Harray[103][186], Harray[104][186], Harray[105][186], Harray[106][186], Harray[107][186], Harray[108][186], Harray[109][186], Harray[110][186], Harray[111][186], Harray[112][186], Harray[113][186], Harray[114][186], Harray[115][186], Harray[116][186], Harray[117][186], Harray[118][186], Harray[119][186], Harray[120][186], Harray[121][186], Harray[122][186], Harray[123][186], Harray[124][186], Harray[125][186], Harray[126][186], Harray[127][186]};
assign h_col_187 = {Harray[0][187], Harray[1][187], Harray[2][187], Harray[3][187], Harray[4][187], Harray[5][187], Harray[6][187], Harray[7][187], Harray[8][187], Harray[9][187], Harray[10][187], Harray[11][187], Harray[12][187], Harray[13][187], Harray[14][187], Harray[15][187], Harray[16][187], Harray[17][187], Harray[18][187], Harray[19][187], Harray[20][187], Harray[21][187], Harray[22][187], Harray[23][187], Harray[24][187], Harray[25][187], Harray[26][187], Harray[27][187], Harray[28][187], Harray[29][187], Harray[30][187], Harray[31][187], Harray[32][187], Harray[33][187], Harray[34][187], Harray[35][187], Harray[36][187], Harray[37][187], Harray[38][187], Harray[39][187], Harray[40][187], Harray[41][187], Harray[42][187], Harray[43][187], Harray[44][187], Harray[45][187], Harray[46][187], Harray[47][187], Harray[48][187], Harray[49][187], Harray[50][187], Harray[51][187], Harray[52][187], Harray[53][187], Harray[54][187], Harray[55][187], Harray[56][187], Harray[57][187], Harray[58][187], Harray[59][187], Harray[60][187], Harray[61][187], Harray[62][187], Harray[63][187], Harray[64][187], Harray[65][187], Harray[66][187], Harray[67][187], Harray[68][187], Harray[69][187], Harray[70][187], Harray[71][187], Harray[72][187], Harray[73][187], Harray[74][187], Harray[75][187], Harray[76][187], Harray[77][187], Harray[78][187], Harray[79][187], Harray[80][187], Harray[81][187], Harray[82][187], Harray[83][187], Harray[84][187], Harray[85][187], Harray[86][187], Harray[87][187], Harray[88][187], Harray[89][187], Harray[90][187], Harray[91][187], Harray[92][187], Harray[93][187], Harray[94][187], Harray[95][187], Harray[96][187], Harray[97][187], Harray[98][187], Harray[99][187], Harray[100][187], Harray[101][187], Harray[102][187], Harray[103][187], Harray[104][187], Harray[105][187], Harray[106][187], Harray[107][187], Harray[108][187], Harray[109][187], Harray[110][187], Harray[111][187], Harray[112][187], Harray[113][187], Harray[114][187], Harray[115][187], Harray[116][187], Harray[117][187], Harray[118][187], Harray[119][187], Harray[120][187], Harray[121][187], Harray[122][187], Harray[123][187], Harray[124][187], Harray[125][187], Harray[126][187], Harray[127][187]};
assign h_col_188 = {Harray[0][188], Harray[1][188], Harray[2][188], Harray[3][188], Harray[4][188], Harray[5][188], Harray[6][188], Harray[7][188], Harray[8][188], Harray[9][188], Harray[10][188], Harray[11][188], Harray[12][188], Harray[13][188], Harray[14][188], Harray[15][188], Harray[16][188], Harray[17][188], Harray[18][188], Harray[19][188], Harray[20][188], Harray[21][188], Harray[22][188], Harray[23][188], Harray[24][188], Harray[25][188], Harray[26][188], Harray[27][188], Harray[28][188], Harray[29][188], Harray[30][188], Harray[31][188], Harray[32][188], Harray[33][188], Harray[34][188], Harray[35][188], Harray[36][188], Harray[37][188], Harray[38][188], Harray[39][188], Harray[40][188], Harray[41][188], Harray[42][188], Harray[43][188], Harray[44][188], Harray[45][188], Harray[46][188], Harray[47][188], Harray[48][188], Harray[49][188], Harray[50][188], Harray[51][188], Harray[52][188], Harray[53][188], Harray[54][188], Harray[55][188], Harray[56][188], Harray[57][188], Harray[58][188], Harray[59][188], Harray[60][188], Harray[61][188], Harray[62][188], Harray[63][188], Harray[64][188], Harray[65][188], Harray[66][188], Harray[67][188], Harray[68][188], Harray[69][188], Harray[70][188], Harray[71][188], Harray[72][188], Harray[73][188], Harray[74][188], Harray[75][188], Harray[76][188], Harray[77][188], Harray[78][188], Harray[79][188], Harray[80][188], Harray[81][188], Harray[82][188], Harray[83][188], Harray[84][188], Harray[85][188], Harray[86][188], Harray[87][188], Harray[88][188], Harray[89][188], Harray[90][188], Harray[91][188], Harray[92][188], Harray[93][188], Harray[94][188], Harray[95][188], Harray[96][188], Harray[97][188], Harray[98][188], Harray[99][188], Harray[100][188], Harray[101][188], Harray[102][188], Harray[103][188], Harray[104][188], Harray[105][188], Harray[106][188], Harray[107][188], Harray[108][188], Harray[109][188], Harray[110][188], Harray[111][188], Harray[112][188], Harray[113][188], Harray[114][188], Harray[115][188], Harray[116][188], Harray[117][188], Harray[118][188], Harray[119][188], Harray[120][188], Harray[121][188], Harray[122][188], Harray[123][188], Harray[124][188], Harray[125][188], Harray[126][188], Harray[127][188]};
assign h_col_189 = {Harray[0][189], Harray[1][189], Harray[2][189], Harray[3][189], Harray[4][189], Harray[5][189], Harray[6][189], Harray[7][189], Harray[8][189], Harray[9][189], Harray[10][189], Harray[11][189], Harray[12][189], Harray[13][189], Harray[14][189], Harray[15][189], Harray[16][189], Harray[17][189], Harray[18][189], Harray[19][189], Harray[20][189], Harray[21][189], Harray[22][189], Harray[23][189], Harray[24][189], Harray[25][189], Harray[26][189], Harray[27][189], Harray[28][189], Harray[29][189], Harray[30][189], Harray[31][189], Harray[32][189], Harray[33][189], Harray[34][189], Harray[35][189], Harray[36][189], Harray[37][189], Harray[38][189], Harray[39][189], Harray[40][189], Harray[41][189], Harray[42][189], Harray[43][189], Harray[44][189], Harray[45][189], Harray[46][189], Harray[47][189], Harray[48][189], Harray[49][189], Harray[50][189], Harray[51][189], Harray[52][189], Harray[53][189], Harray[54][189], Harray[55][189], Harray[56][189], Harray[57][189], Harray[58][189], Harray[59][189], Harray[60][189], Harray[61][189], Harray[62][189], Harray[63][189], Harray[64][189], Harray[65][189], Harray[66][189], Harray[67][189], Harray[68][189], Harray[69][189], Harray[70][189], Harray[71][189], Harray[72][189], Harray[73][189], Harray[74][189], Harray[75][189], Harray[76][189], Harray[77][189], Harray[78][189], Harray[79][189], Harray[80][189], Harray[81][189], Harray[82][189], Harray[83][189], Harray[84][189], Harray[85][189], Harray[86][189], Harray[87][189], Harray[88][189], Harray[89][189], Harray[90][189], Harray[91][189], Harray[92][189], Harray[93][189], Harray[94][189], Harray[95][189], Harray[96][189], Harray[97][189], Harray[98][189], Harray[99][189], Harray[100][189], Harray[101][189], Harray[102][189], Harray[103][189], Harray[104][189], Harray[105][189], Harray[106][189], Harray[107][189], Harray[108][189], Harray[109][189], Harray[110][189], Harray[111][189], Harray[112][189], Harray[113][189], Harray[114][189], Harray[115][189], Harray[116][189], Harray[117][189], Harray[118][189], Harray[119][189], Harray[120][189], Harray[121][189], Harray[122][189], Harray[123][189], Harray[124][189], Harray[125][189], Harray[126][189], Harray[127][189]};
assign h_col_190 = {Harray[0][190], Harray[1][190], Harray[2][190], Harray[3][190], Harray[4][190], Harray[5][190], Harray[6][190], Harray[7][190], Harray[8][190], Harray[9][190], Harray[10][190], Harray[11][190], Harray[12][190], Harray[13][190], Harray[14][190], Harray[15][190], Harray[16][190], Harray[17][190], Harray[18][190], Harray[19][190], Harray[20][190], Harray[21][190], Harray[22][190], Harray[23][190], Harray[24][190], Harray[25][190], Harray[26][190], Harray[27][190], Harray[28][190], Harray[29][190], Harray[30][190], Harray[31][190], Harray[32][190], Harray[33][190], Harray[34][190], Harray[35][190], Harray[36][190], Harray[37][190], Harray[38][190], Harray[39][190], Harray[40][190], Harray[41][190], Harray[42][190], Harray[43][190], Harray[44][190], Harray[45][190], Harray[46][190], Harray[47][190], Harray[48][190], Harray[49][190], Harray[50][190], Harray[51][190], Harray[52][190], Harray[53][190], Harray[54][190], Harray[55][190], Harray[56][190], Harray[57][190], Harray[58][190], Harray[59][190], Harray[60][190], Harray[61][190], Harray[62][190], Harray[63][190], Harray[64][190], Harray[65][190], Harray[66][190], Harray[67][190], Harray[68][190], Harray[69][190], Harray[70][190], Harray[71][190], Harray[72][190], Harray[73][190], Harray[74][190], Harray[75][190], Harray[76][190], Harray[77][190], Harray[78][190], Harray[79][190], Harray[80][190], Harray[81][190], Harray[82][190], Harray[83][190], Harray[84][190], Harray[85][190], Harray[86][190], Harray[87][190], Harray[88][190], Harray[89][190], Harray[90][190], Harray[91][190], Harray[92][190], Harray[93][190], Harray[94][190], Harray[95][190], Harray[96][190], Harray[97][190], Harray[98][190], Harray[99][190], Harray[100][190], Harray[101][190], Harray[102][190], Harray[103][190], Harray[104][190], Harray[105][190], Harray[106][190], Harray[107][190], Harray[108][190], Harray[109][190], Harray[110][190], Harray[111][190], Harray[112][190], Harray[113][190], Harray[114][190], Harray[115][190], Harray[116][190], Harray[117][190], Harray[118][190], Harray[119][190], Harray[120][190], Harray[121][190], Harray[122][190], Harray[123][190], Harray[124][190], Harray[125][190], Harray[126][190], Harray[127][190]};
assign h_col_191 = {Harray[0][191], Harray[1][191], Harray[2][191], Harray[3][191], Harray[4][191], Harray[5][191], Harray[6][191], Harray[7][191], Harray[8][191], Harray[9][191], Harray[10][191], Harray[11][191], Harray[12][191], Harray[13][191], Harray[14][191], Harray[15][191], Harray[16][191], Harray[17][191], Harray[18][191], Harray[19][191], Harray[20][191], Harray[21][191], Harray[22][191], Harray[23][191], Harray[24][191], Harray[25][191], Harray[26][191], Harray[27][191], Harray[28][191], Harray[29][191], Harray[30][191], Harray[31][191], Harray[32][191], Harray[33][191], Harray[34][191], Harray[35][191], Harray[36][191], Harray[37][191], Harray[38][191], Harray[39][191], Harray[40][191], Harray[41][191], Harray[42][191], Harray[43][191], Harray[44][191], Harray[45][191], Harray[46][191], Harray[47][191], Harray[48][191], Harray[49][191], Harray[50][191], Harray[51][191], Harray[52][191], Harray[53][191], Harray[54][191], Harray[55][191], Harray[56][191], Harray[57][191], Harray[58][191], Harray[59][191], Harray[60][191], Harray[61][191], Harray[62][191], Harray[63][191], Harray[64][191], Harray[65][191], Harray[66][191], Harray[67][191], Harray[68][191], Harray[69][191], Harray[70][191], Harray[71][191], Harray[72][191], Harray[73][191], Harray[74][191], Harray[75][191], Harray[76][191], Harray[77][191], Harray[78][191], Harray[79][191], Harray[80][191], Harray[81][191], Harray[82][191], Harray[83][191], Harray[84][191], Harray[85][191], Harray[86][191], Harray[87][191], Harray[88][191], Harray[89][191], Harray[90][191], Harray[91][191], Harray[92][191], Harray[93][191], Harray[94][191], Harray[95][191], Harray[96][191], Harray[97][191], Harray[98][191], Harray[99][191], Harray[100][191], Harray[101][191], Harray[102][191], Harray[103][191], Harray[104][191], Harray[105][191], Harray[106][191], Harray[107][191], Harray[108][191], Harray[109][191], Harray[110][191], Harray[111][191], Harray[112][191], Harray[113][191], Harray[114][191], Harray[115][191], Harray[116][191], Harray[117][191], Harray[118][191], Harray[119][191], Harray[120][191], Harray[121][191], Harray[122][191], Harray[123][191], Harray[124][191], Harray[125][191], Harray[126][191], Harray[127][191]};
assign h_col_192 = {Harray[0][192], Harray[1][192], Harray[2][192], Harray[3][192], Harray[4][192], Harray[5][192], Harray[6][192], Harray[7][192], Harray[8][192], Harray[9][192], Harray[10][192], Harray[11][192], Harray[12][192], Harray[13][192], Harray[14][192], Harray[15][192], Harray[16][192], Harray[17][192], Harray[18][192], Harray[19][192], Harray[20][192], Harray[21][192], Harray[22][192], Harray[23][192], Harray[24][192], Harray[25][192], Harray[26][192], Harray[27][192], Harray[28][192], Harray[29][192], Harray[30][192], Harray[31][192], Harray[32][192], Harray[33][192], Harray[34][192], Harray[35][192], Harray[36][192], Harray[37][192], Harray[38][192], Harray[39][192], Harray[40][192], Harray[41][192], Harray[42][192], Harray[43][192], Harray[44][192], Harray[45][192], Harray[46][192], Harray[47][192], Harray[48][192], Harray[49][192], Harray[50][192], Harray[51][192], Harray[52][192], Harray[53][192], Harray[54][192], Harray[55][192], Harray[56][192], Harray[57][192], Harray[58][192], Harray[59][192], Harray[60][192], Harray[61][192], Harray[62][192], Harray[63][192], Harray[64][192], Harray[65][192], Harray[66][192], Harray[67][192], Harray[68][192], Harray[69][192], Harray[70][192], Harray[71][192], Harray[72][192], Harray[73][192], Harray[74][192], Harray[75][192], Harray[76][192], Harray[77][192], Harray[78][192], Harray[79][192], Harray[80][192], Harray[81][192], Harray[82][192], Harray[83][192], Harray[84][192], Harray[85][192], Harray[86][192], Harray[87][192], Harray[88][192], Harray[89][192], Harray[90][192], Harray[91][192], Harray[92][192], Harray[93][192], Harray[94][192], Harray[95][192], Harray[96][192], Harray[97][192], Harray[98][192], Harray[99][192], Harray[100][192], Harray[101][192], Harray[102][192], Harray[103][192], Harray[104][192], Harray[105][192], Harray[106][192], Harray[107][192], Harray[108][192], Harray[109][192], Harray[110][192], Harray[111][192], Harray[112][192], Harray[113][192], Harray[114][192], Harray[115][192], Harray[116][192], Harray[117][192], Harray[118][192], Harray[119][192], Harray[120][192], Harray[121][192], Harray[122][192], Harray[123][192], Harray[124][192], Harray[125][192], Harray[126][192], Harray[127][192]};
assign h_col_193 = {Harray[0][193], Harray[1][193], Harray[2][193], Harray[3][193], Harray[4][193], Harray[5][193], Harray[6][193], Harray[7][193], Harray[8][193], Harray[9][193], Harray[10][193], Harray[11][193], Harray[12][193], Harray[13][193], Harray[14][193], Harray[15][193], Harray[16][193], Harray[17][193], Harray[18][193], Harray[19][193], Harray[20][193], Harray[21][193], Harray[22][193], Harray[23][193], Harray[24][193], Harray[25][193], Harray[26][193], Harray[27][193], Harray[28][193], Harray[29][193], Harray[30][193], Harray[31][193], Harray[32][193], Harray[33][193], Harray[34][193], Harray[35][193], Harray[36][193], Harray[37][193], Harray[38][193], Harray[39][193], Harray[40][193], Harray[41][193], Harray[42][193], Harray[43][193], Harray[44][193], Harray[45][193], Harray[46][193], Harray[47][193], Harray[48][193], Harray[49][193], Harray[50][193], Harray[51][193], Harray[52][193], Harray[53][193], Harray[54][193], Harray[55][193], Harray[56][193], Harray[57][193], Harray[58][193], Harray[59][193], Harray[60][193], Harray[61][193], Harray[62][193], Harray[63][193], Harray[64][193], Harray[65][193], Harray[66][193], Harray[67][193], Harray[68][193], Harray[69][193], Harray[70][193], Harray[71][193], Harray[72][193], Harray[73][193], Harray[74][193], Harray[75][193], Harray[76][193], Harray[77][193], Harray[78][193], Harray[79][193], Harray[80][193], Harray[81][193], Harray[82][193], Harray[83][193], Harray[84][193], Harray[85][193], Harray[86][193], Harray[87][193], Harray[88][193], Harray[89][193], Harray[90][193], Harray[91][193], Harray[92][193], Harray[93][193], Harray[94][193], Harray[95][193], Harray[96][193], Harray[97][193], Harray[98][193], Harray[99][193], Harray[100][193], Harray[101][193], Harray[102][193], Harray[103][193], Harray[104][193], Harray[105][193], Harray[106][193], Harray[107][193], Harray[108][193], Harray[109][193], Harray[110][193], Harray[111][193], Harray[112][193], Harray[113][193], Harray[114][193], Harray[115][193], Harray[116][193], Harray[117][193], Harray[118][193], Harray[119][193], Harray[120][193], Harray[121][193], Harray[122][193], Harray[123][193], Harray[124][193], Harray[125][193], Harray[126][193], Harray[127][193]};
assign h_col_194 = {Harray[0][194], Harray[1][194], Harray[2][194], Harray[3][194], Harray[4][194], Harray[5][194], Harray[6][194], Harray[7][194], Harray[8][194], Harray[9][194], Harray[10][194], Harray[11][194], Harray[12][194], Harray[13][194], Harray[14][194], Harray[15][194], Harray[16][194], Harray[17][194], Harray[18][194], Harray[19][194], Harray[20][194], Harray[21][194], Harray[22][194], Harray[23][194], Harray[24][194], Harray[25][194], Harray[26][194], Harray[27][194], Harray[28][194], Harray[29][194], Harray[30][194], Harray[31][194], Harray[32][194], Harray[33][194], Harray[34][194], Harray[35][194], Harray[36][194], Harray[37][194], Harray[38][194], Harray[39][194], Harray[40][194], Harray[41][194], Harray[42][194], Harray[43][194], Harray[44][194], Harray[45][194], Harray[46][194], Harray[47][194], Harray[48][194], Harray[49][194], Harray[50][194], Harray[51][194], Harray[52][194], Harray[53][194], Harray[54][194], Harray[55][194], Harray[56][194], Harray[57][194], Harray[58][194], Harray[59][194], Harray[60][194], Harray[61][194], Harray[62][194], Harray[63][194], Harray[64][194], Harray[65][194], Harray[66][194], Harray[67][194], Harray[68][194], Harray[69][194], Harray[70][194], Harray[71][194], Harray[72][194], Harray[73][194], Harray[74][194], Harray[75][194], Harray[76][194], Harray[77][194], Harray[78][194], Harray[79][194], Harray[80][194], Harray[81][194], Harray[82][194], Harray[83][194], Harray[84][194], Harray[85][194], Harray[86][194], Harray[87][194], Harray[88][194], Harray[89][194], Harray[90][194], Harray[91][194], Harray[92][194], Harray[93][194], Harray[94][194], Harray[95][194], Harray[96][194], Harray[97][194], Harray[98][194], Harray[99][194], Harray[100][194], Harray[101][194], Harray[102][194], Harray[103][194], Harray[104][194], Harray[105][194], Harray[106][194], Harray[107][194], Harray[108][194], Harray[109][194], Harray[110][194], Harray[111][194], Harray[112][194], Harray[113][194], Harray[114][194], Harray[115][194], Harray[116][194], Harray[117][194], Harray[118][194], Harray[119][194], Harray[120][194], Harray[121][194], Harray[122][194], Harray[123][194], Harray[124][194], Harray[125][194], Harray[126][194], Harray[127][194]};
assign h_col_195 = {Harray[0][195], Harray[1][195], Harray[2][195], Harray[3][195], Harray[4][195], Harray[5][195], Harray[6][195], Harray[7][195], Harray[8][195], Harray[9][195], Harray[10][195], Harray[11][195], Harray[12][195], Harray[13][195], Harray[14][195], Harray[15][195], Harray[16][195], Harray[17][195], Harray[18][195], Harray[19][195], Harray[20][195], Harray[21][195], Harray[22][195], Harray[23][195], Harray[24][195], Harray[25][195], Harray[26][195], Harray[27][195], Harray[28][195], Harray[29][195], Harray[30][195], Harray[31][195], Harray[32][195], Harray[33][195], Harray[34][195], Harray[35][195], Harray[36][195], Harray[37][195], Harray[38][195], Harray[39][195], Harray[40][195], Harray[41][195], Harray[42][195], Harray[43][195], Harray[44][195], Harray[45][195], Harray[46][195], Harray[47][195], Harray[48][195], Harray[49][195], Harray[50][195], Harray[51][195], Harray[52][195], Harray[53][195], Harray[54][195], Harray[55][195], Harray[56][195], Harray[57][195], Harray[58][195], Harray[59][195], Harray[60][195], Harray[61][195], Harray[62][195], Harray[63][195], Harray[64][195], Harray[65][195], Harray[66][195], Harray[67][195], Harray[68][195], Harray[69][195], Harray[70][195], Harray[71][195], Harray[72][195], Harray[73][195], Harray[74][195], Harray[75][195], Harray[76][195], Harray[77][195], Harray[78][195], Harray[79][195], Harray[80][195], Harray[81][195], Harray[82][195], Harray[83][195], Harray[84][195], Harray[85][195], Harray[86][195], Harray[87][195], Harray[88][195], Harray[89][195], Harray[90][195], Harray[91][195], Harray[92][195], Harray[93][195], Harray[94][195], Harray[95][195], Harray[96][195], Harray[97][195], Harray[98][195], Harray[99][195], Harray[100][195], Harray[101][195], Harray[102][195], Harray[103][195], Harray[104][195], Harray[105][195], Harray[106][195], Harray[107][195], Harray[108][195], Harray[109][195], Harray[110][195], Harray[111][195], Harray[112][195], Harray[113][195], Harray[114][195], Harray[115][195], Harray[116][195], Harray[117][195], Harray[118][195], Harray[119][195], Harray[120][195], Harray[121][195], Harray[122][195], Harray[123][195], Harray[124][195], Harray[125][195], Harray[126][195], Harray[127][195]};
assign h_col_196 = {Harray[0][196], Harray[1][196], Harray[2][196], Harray[3][196], Harray[4][196], Harray[5][196], Harray[6][196], Harray[7][196], Harray[8][196], Harray[9][196], Harray[10][196], Harray[11][196], Harray[12][196], Harray[13][196], Harray[14][196], Harray[15][196], Harray[16][196], Harray[17][196], Harray[18][196], Harray[19][196], Harray[20][196], Harray[21][196], Harray[22][196], Harray[23][196], Harray[24][196], Harray[25][196], Harray[26][196], Harray[27][196], Harray[28][196], Harray[29][196], Harray[30][196], Harray[31][196], Harray[32][196], Harray[33][196], Harray[34][196], Harray[35][196], Harray[36][196], Harray[37][196], Harray[38][196], Harray[39][196], Harray[40][196], Harray[41][196], Harray[42][196], Harray[43][196], Harray[44][196], Harray[45][196], Harray[46][196], Harray[47][196], Harray[48][196], Harray[49][196], Harray[50][196], Harray[51][196], Harray[52][196], Harray[53][196], Harray[54][196], Harray[55][196], Harray[56][196], Harray[57][196], Harray[58][196], Harray[59][196], Harray[60][196], Harray[61][196], Harray[62][196], Harray[63][196], Harray[64][196], Harray[65][196], Harray[66][196], Harray[67][196], Harray[68][196], Harray[69][196], Harray[70][196], Harray[71][196], Harray[72][196], Harray[73][196], Harray[74][196], Harray[75][196], Harray[76][196], Harray[77][196], Harray[78][196], Harray[79][196], Harray[80][196], Harray[81][196], Harray[82][196], Harray[83][196], Harray[84][196], Harray[85][196], Harray[86][196], Harray[87][196], Harray[88][196], Harray[89][196], Harray[90][196], Harray[91][196], Harray[92][196], Harray[93][196], Harray[94][196], Harray[95][196], Harray[96][196], Harray[97][196], Harray[98][196], Harray[99][196], Harray[100][196], Harray[101][196], Harray[102][196], Harray[103][196], Harray[104][196], Harray[105][196], Harray[106][196], Harray[107][196], Harray[108][196], Harray[109][196], Harray[110][196], Harray[111][196], Harray[112][196], Harray[113][196], Harray[114][196], Harray[115][196], Harray[116][196], Harray[117][196], Harray[118][196], Harray[119][196], Harray[120][196], Harray[121][196], Harray[122][196], Harray[123][196], Harray[124][196], Harray[125][196], Harray[126][196], Harray[127][196]};
assign h_col_197 = {Harray[0][197], Harray[1][197], Harray[2][197], Harray[3][197], Harray[4][197], Harray[5][197], Harray[6][197], Harray[7][197], Harray[8][197], Harray[9][197], Harray[10][197], Harray[11][197], Harray[12][197], Harray[13][197], Harray[14][197], Harray[15][197], Harray[16][197], Harray[17][197], Harray[18][197], Harray[19][197], Harray[20][197], Harray[21][197], Harray[22][197], Harray[23][197], Harray[24][197], Harray[25][197], Harray[26][197], Harray[27][197], Harray[28][197], Harray[29][197], Harray[30][197], Harray[31][197], Harray[32][197], Harray[33][197], Harray[34][197], Harray[35][197], Harray[36][197], Harray[37][197], Harray[38][197], Harray[39][197], Harray[40][197], Harray[41][197], Harray[42][197], Harray[43][197], Harray[44][197], Harray[45][197], Harray[46][197], Harray[47][197], Harray[48][197], Harray[49][197], Harray[50][197], Harray[51][197], Harray[52][197], Harray[53][197], Harray[54][197], Harray[55][197], Harray[56][197], Harray[57][197], Harray[58][197], Harray[59][197], Harray[60][197], Harray[61][197], Harray[62][197], Harray[63][197], Harray[64][197], Harray[65][197], Harray[66][197], Harray[67][197], Harray[68][197], Harray[69][197], Harray[70][197], Harray[71][197], Harray[72][197], Harray[73][197], Harray[74][197], Harray[75][197], Harray[76][197], Harray[77][197], Harray[78][197], Harray[79][197], Harray[80][197], Harray[81][197], Harray[82][197], Harray[83][197], Harray[84][197], Harray[85][197], Harray[86][197], Harray[87][197], Harray[88][197], Harray[89][197], Harray[90][197], Harray[91][197], Harray[92][197], Harray[93][197], Harray[94][197], Harray[95][197], Harray[96][197], Harray[97][197], Harray[98][197], Harray[99][197], Harray[100][197], Harray[101][197], Harray[102][197], Harray[103][197], Harray[104][197], Harray[105][197], Harray[106][197], Harray[107][197], Harray[108][197], Harray[109][197], Harray[110][197], Harray[111][197], Harray[112][197], Harray[113][197], Harray[114][197], Harray[115][197], Harray[116][197], Harray[117][197], Harray[118][197], Harray[119][197], Harray[120][197], Harray[121][197], Harray[122][197], Harray[123][197], Harray[124][197], Harray[125][197], Harray[126][197], Harray[127][197]};
assign h_col_198 = {Harray[0][198], Harray[1][198], Harray[2][198], Harray[3][198], Harray[4][198], Harray[5][198], Harray[6][198], Harray[7][198], Harray[8][198], Harray[9][198], Harray[10][198], Harray[11][198], Harray[12][198], Harray[13][198], Harray[14][198], Harray[15][198], Harray[16][198], Harray[17][198], Harray[18][198], Harray[19][198], Harray[20][198], Harray[21][198], Harray[22][198], Harray[23][198], Harray[24][198], Harray[25][198], Harray[26][198], Harray[27][198], Harray[28][198], Harray[29][198], Harray[30][198], Harray[31][198], Harray[32][198], Harray[33][198], Harray[34][198], Harray[35][198], Harray[36][198], Harray[37][198], Harray[38][198], Harray[39][198], Harray[40][198], Harray[41][198], Harray[42][198], Harray[43][198], Harray[44][198], Harray[45][198], Harray[46][198], Harray[47][198], Harray[48][198], Harray[49][198], Harray[50][198], Harray[51][198], Harray[52][198], Harray[53][198], Harray[54][198], Harray[55][198], Harray[56][198], Harray[57][198], Harray[58][198], Harray[59][198], Harray[60][198], Harray[61][198], Harray[62][198], Harray[63][198], Harray[64][198], Harray[65][198], Harray[66][198], Harray[67][198], Harray[68][198], Harray[69][198], Harray[70][198], Harray[71][198], Harray[72][198], Harray[73][198], Harray[74][198], Harray[75][198], Harray[76][198], Harray[77][198], Harray[78][198], Harray[79][198], Harray[80][198], Harray[81][198], Harray[82][198], Harray[83][198], Harray[84][198], Harray[85][198], Harray[86][198], Harray[87][198], Harray[88][198], Harray[89][198], Harray[90][198], Harray[91][198], Harray[92][198], Harray[93][198], Harray[94][198], Harray[95][198], Harray[96][198], Harray[97][198], Harray[98][198], Harray[99][198], Harray[100][198], Harray[101][198], Harray[102][198], Harray[103][198], Harray[104][198], Harray[105][198], Harray[106][198], Harray[107][198], Harray[108][198], Harray[109][198], Harray[110][198], Harray[111][198], Harray[112][198], Harray[113][198], Harray[114][198], Harray[115][198], Harray[116][198], Harray[117][198], Harray[118][198], Harray[119][198], Harray[120][198], Harray[121][198], Harray[122][198], Harray[123][198], Harray[124][198], Harray[125][198], Harray[126][198], Harray[127][198]};
assign h_col_199 = {Harray[0][199], Harray[1][199], Harray[2][199], Harray[3][199], Harray[4][199], Harray[5][199], Harray[6][199], Harray[7][199], Harray[8][199], Harray[9][199], Harray[10][199], Harray[11][199], Harray[12][199], Harray[13][199], Harray[14][199], Harray[15][199], Harray[16][199], Harray[17][199], Harray[18][199], Harray[19][199], Harray[20][199], Harray[21][199], Harray[22][199], Harray[23][199], Harray[24][199], Harray[25][199], Harray[26][199], Harray[27][199], Harray[28][199], Harray[29][199], Harray[30][199], Harray[31][199], Harray[32][199], Harray[33][199], Harray[34][199], Harray[35][199], Harray[36][199], Harray[37][199], Harray[38][199], Harray[39][199], Harray[40][199], Harray[41][199], Harray[42][199], Harray[43][199], Harray[44][199], Harray[45][199], Harray[46][199], Harray[47][199], Harray[48][199], Harray[49][199], Harray[50][199], Harray[51][199], Harray[52][199], Harray[53][199], Harray[54][199], Harray[55][199], Harray[56][199], Harray[57][199], Harray[58][199], Harray[59][199], Harray[60][199], Harray[61][199], Harray[62][199], Harray[63][199], Harray[64][199], Harray[65][199], Harray[66][199], Harray[67][199], Harray[68][199], Harray[69][199], Harray[70][199], Harray[71][199], Harray[72][199], Harray[73][199], Harray[74][199], Harray[75][199], Harray[76][199], Harray[77][199], Harray[78][199], Harray[79][199], Harray[80][199], Harray[81][199], Harray[82][199], Harray[83][199], Harray[84][199], Harray[85][199], Harray[86][199], Harray[87][199], Harray[88][199], Harray[89][199], Harray[90][199], Harray[91][199], Harray[92][199], Harray[93][199], Harray[94][199], Harray[95][199], Harray[96][199], Harray[97][199], Harray[98][199], Harray[99][199], Harray[100][199], Harray[101][199], Harray[102][199], Harray[103][199], Harray[104][199], Harray[105][199], Harray[106][199], Harray[107][199], Harray[108][199], Harray[109][199], Harray[110][199], Harray[111][199], Harray[112][199], Harray[113][199], Harray[114][199], Harray[115][199], Harray[116][199], Harray[117][199], Harray[118][199], Harray[119][199], Harray[120][199], Harray[121][199], Harray[122][199], Harray[123][199], Harray[124][199], Harray[125][199], Harray[126][199], Harray[127][199]};
assign h_col_200 = {Harray[0][200], Harray[1][200], Harray[2][200], Harray[3][200], Harray[4][200], Harray[5][200], Harray[6][200], Harray[7][200], Harray[8][200], Harray[9][200], Harray[10][200], Harray[11][200], Harray[12][200], Harray[13][200], Harray[14][200], Harray[15][200], Harray[16][200], Harray[17][200], Harray[18][200], Harray[19][200], Harray[20][200], Harray[21][200], Harray[22][200], Harray[23][200], Harray[24][200], Harray[25][200], Harray[26][200], Harray[27][200], Harray[28][200], Harray[29][200], Harray[30][200], Harray[31][200], Harray[32][200], Harray[33][200], Harray[34][200], Harray[35][200], Harray[36][200], Harray[37][200], Harray[38][200], Harray[39][200], Harray[40][200], Harray[41][200], Harray[42][200], Harray[43][200], Harray[44][200], Harray[45][200], Harray[46][200], Harray[47][200], Harray[48][200], Harray[49][200], Harray[50][200], Harray[51][200], Harray[52][200], Harray[53][200], Harray[54][200], Harray[55][200], Harray[56][200], Harray[57][200], Harray[58][200], Harray[59][200], Harray[60][200], Harray[61][200], Harray[62][200], Harray[63][200], Harray[64][200], Harray[65][200], Harray[66][200], Harray[67][200], Harray[68][200], Harray[69][200], Harray[70][200], Harray[71][200], Harray[72][200], Harray[73][200], Harray[74][200], Harray[75][200], Harray[76][200], Harray[77][200], Harray[78][200], Harray[79][200], Harray[80][200], Harray[81][200], Harray[82][200], Harray[83][200], Harray[84][200], Harray[85][200], Harray[86][200], Harray[87][200], Harray[88][200], Harray[89][200], Harray[90][200], Harray[91][200], Harray[92][200], Harray[93][200], Harray[94][200], Harray[95][200], Harray[96][200], Harray[97][200], Harray[98][200], Harray[99][200], Harray[100][200], Harray[101][200], Harray[102][200], Harray[103][200], Harray[104][200], Harray[105][200], Harray[106][200], Harray[107][200], Harray[108][200], Harray[109][200], Harray[110][200], Harray[111][200], Harray[112][200], Harray[113][200], Harray[114][200], Harray[115][200], Harray[116][200], Harray[117][200], Harray[118][200], Harray[119][200], Harray[120][200], Harray[121][200], Harray[122][200], Harray[123][200], Harray[124][200], Harray[125][200], Harray[126][200], Harray[127][200]};
assign h_col_201 = {Harray[0][201], Harray[1][201], Harray[2][201], Harray[3][201], Harray[4][201], Harray[5][201], Harray[6][201], Harray[7][201], Harray[8][201], Harray[9][201], Harray[10][201], Harray[11][201], Harray[12][201], Harray[13][201], Harray[14][201], Harray[15][201], Harray[16][201], Harray[17][201], Harray[18][201], Harray[19][201], Harray[20][201], Harray[21][201], Harray[22][201], Harray[23][201], Harray[24][201], Harray[25][201], Harray[26][201], Harray[27][201], Harray[28][201], Harray[29][201], Harray[30][201], Harray[31][201], Harray[32][201], Harray[33][201], Harray[34][201], Harray[35][201], Harray[36][201], Harray[37][201], Harray[38][201], Harray[39][201], Harray[40][201], Harray[41][201], Harray[42][201], Harray[43][201], Harray[44][201], Harray[45][201], Harray[46][201], Harray[47][201], Harray[48][201], Harray[49][201], Harray[50][201], Harray[51][201], Harray[52][201], Harray[53][201], Harray[54][201], Harray[55][201], Harray[56][201], Harray[57][201], Harray[58][201], Harray[59][201], Harray[60][201], Harray[61][201], Harray[62][201], Harray[63][201], Harray[64][201], Harray[65][201], Harray[66][201], Harray[67][201], Harray[68][201], Harray[69][201], Harray[70][201], Harray[71][201], Harray[72][201], Harray[73][201], Harray[74][201], Harray[75][201], Harray[76][201], Harray[77][201], Harray[78][201], Harray[79][201], Harray[80][201], Harray[81][201], Harray[82][201], Harray[83][201], Harray[84][201], Harray[85][201], Harray[86][201], Harray[87][201], Harray[88][201], Harray[89][201], Harray[90][201], Harray[91][201], Harray[92][201], Harray[93][201], Harray[94][201], Harray[95][201], Harray[96][201], Harray[97][201], Harray[98][201], Harray[99][201], Harray[100][201], Harray[101][201], Harray[102][201], Harray[103][201], Harray[104][201], Harray[105][201], Harray[106][201], Harray[107][201], Harray[108][201], Harray[109][201], Harray[110][201], Harray[111][201], Harray[112][201], Harray[113][201], Harray[114][201], Harray[115][201], Harray[116][201], Harray[117][201], Harray[118][201], Harray[119][201], Harray[120][201], Harray[121][201], Harray[122][201], Harray[123][201], Harray[124][201], Harray[125][201], Harray[126][201], Harray[127][201]};
assign h_col_202 = {Harray[0][202], Harray[1][202], Harray[2][202], Harray[3][202], Harray[4][202], Harray[5][202], Harray[6][202], Harray[7][202], Harray[8][202], Harray[9][202], Harray[10][202], Harray[11][202], Harray[12][202], Harray[13][202], Harray[14][202], Harray[15][202], Harray[16][202], Harray[17][202], Harray[18][202], Harray[19][202], Harray[20][202], Harray[21][202], Harray[22][202], Harray[23][202], Harray[24][202], Harray[25][202], Harray[26][202], Harray[27][202], Harray[28][202], Harray[29][202], Harray[30][202], Harray[31][202], Harray[32][202], Harray[33][202], Harray[34][202], Harray[35][202], Harray[36][202], Harray[37][202], Harray[38][202], Harray[39][202], Harray[40][202], Harray[41][202], Harray[42][202], Harray[43][202], Harray[44][202], Harray[45][202], Harray[46][202], Harray[47][202], Harray[48][202], Harray[49][202], Harray[50][202], Harray[51][202], Harray[52][202], Harray[53][202], Harray[54][202], Harray[55][202], Harray[56][202], Harray[57][202], Harray[58][202], Harray[59][202], Harray[60][202], Harray[61][202], Harray[62][202], Harray[63][202], Harray[64][202], Harray[65][202], Harray[66][202], Harray[67][202], Harray[68][202], Harray[69][202], Harray[70][202], Harray[71][202], Harray[72][202], Harray[73][202], Harray[74][202], Harray[75][202], Harray[76][202], Harray[77][202], Harray[78][202], Harray[79][202], Harray[80][202], Harray[81][202], Harray[82][202], Harray[83][202], Harray[84][202], Harray[85][202], Harray[86][202], Harray[87][202], Harray[88][202], Harray[89][202], Harray[90][202], Harray[91][202], Harray[92][202], Harray[93][202], Harray[94][202], Harray[95][202], Harray[96][202], Harray[97][202], Harray[98][202], Harray[99][202], Harray[100][202], Harray[101][202], Harray[102][202], Harray[103][202], Harray[104][202], Harray[105][202], Harray[106][202], Harray[107][202], Harray[108][202], Harray[109][202], Harray[110][202], Harray[111][202], Harray[112][202], Harray[113][202], Harray[114][202], Harray[115][202], Harray[116][202], Harray[117][202], Harray[118][202], Harray[119][202], Harray[120][202], Harray[121][202], Harray[122][202], Harray[123][202], Harray[124][202], Harray[125][202], Harray[126][202], Harray[127][202]};
assign h_col_203 = {Harray[0][203], Harray[1][203], Harray[2][203], Harray[3][203], Harray[4][203], Harray[5][203], Harray[6][203], Harray[7][203], Harray[8][203], Harray[9][203], Harray[10][203], Harray[11][203], Harray[12][203], Harray[13][203], Harray[14][203], Harray[15][203], Harray[16][203], Harray[17][203], Harray[18][203], Harray[19][203], Harray[20][203], Harray[21][203], Harray[22][203], Harray[23][203], Harray[24][203], Harray[25][203], Harray[26][203], Harray[27][203], Harray[28][203], Harray[29][203], Harray[30][203], Harray[31][203], Harray[32][203], Harray[33][203], Harray[34][203], Harray[35][203], Harray[36][203], Harray[37][203], Harray[38][203], Harray[39][203], Harray[40][203], Harray[41][203], Harray[42][203], Harray[43][203], Harray[44][203], Harray[45][203], Harray[46][203], Harray[47][203], Harray[48][203], Harray[49][203], Harray[50][203], Harray[51][203], Harray[52][203], Harray[53][203], Harray[54][203], Harray[55][203], Harray[56][203], Harray[57][203], Harray[58][203], Harray[59][203], Harray[60][203], Harray[61][203], Harray[62][203], Harray[63][203], Harray[64][203], Harray[65][203], Harray[66][203], Harray[67][203], Harray[68][203], Harray[69][203], Harray[70][203], Harray[71][203], Harray[72][203], Harray[73][203], Harray[74][203], Harray[75][203], Harray[76][203], Harray[77][203], Harray[78][203], Harray[79][203], Harray[80][203], Harray[81][203], Harray[82][203], Harray[83][203], Harray[84][203], Harray[85][203], Harray[86][203], Harray[87][203], Harray[88][203], Harray[89][203], Harray[90][203], Harray[91][203], Harray[92][203], Harray[93][203], Harray[94][203], Harray[95][203], Harray[96][203], Harray[97][203], Harray[98][203], Harray[99][203], Harray[100][203], Harray[101][203], Harray[102][203], Harray[103][203], Harray[104][203], Harray[105][203], Harray[106][203], Harray[107][203], Harray[108][203], Harray[109][203], Harray[110][203], Harray[111][203], Harray[112][203], Harray[113][203], Harray[114][203], Harray[115][203], Harray[116][203], Harray[117][203], Harray[118][203], Harray[119][203], Harray[120][203], Harray[121][203], Harray[122][203], Harray[123][203], Harray[124][203], Harray[125][203], Harray[126][203], Harray[127][203]};
assign h_col_204 = {Harray[0][204], Harray[1][204], Harray[2][204], Harray[3][204], Harray[4][204], Harray[5][204], Harray[6][204], Harray[7][204], Harray[8][204], Harray[9][204], Harray[10][204], Harray[11][204], Harray[12][204], Harray[13][204], Harray[14][204], Harray[15][204], Harray[16][204], Harray[17][204], Harray[18][204], Harray[19][204], Harray[20][204], Harray[21][204], Harray[22][204], Harray[23][204], Harray[24][204], Harray[25][204], Harray[26][204], Harray[27][204], Harray[28][204], Harray[29][204], Harray[30][204], Harray[31][204], Harray[32][204], Harray[33][204], Harray[34][204], Harray[35][204], Harray[36][204], Harray[37][204], Harray[38][204], Harray[39][204], Harray[40][204], Harray[41][204], Harray[42][204], Harray[43][204], Harray[44][204], Harray[45][204], Harray[46][204], Harray[47][204], Harray[48][204], Harray[49][204], Harray[50][204], Harray[51][204], Harray[52][204], Harray[53][204], Harray[54][204], Harray[55][204], Harray[56][204], Harray[57][204], Harray[58][204], Harray[59][204], Harray[60][204], Harray[61][204], Harray[62][204], Harray[63][204], Harray[64][204], Harray[65][204], Harray[66][204], Harray[67][204], Harray[68][204], Harray[69][204], Harray[70][204], Harray[71][204], Harray[72][204], Harray[73][204], Harray[74][204], Harray[75][204], Harray[76][204], Harray[77][204], Harray[78][204], Harray[79][204], Harray[80][204], Harray[81][204], Harray[82][204], Harray[83][204], Harray[84][204], Harray[85][204], Harray[86][204], Harray[87][204], Harray[88][204], Harray[89][204], Harray[90][204], Harray[91][204], Harray[92][204], Harray[93][204], Harray[94][204], Harray[95][204], Harray[96][204], Harray[97][204], Harray[98][204], Harray[99][204], Harray[100][204], Harray[101][204], Harray[102][204], Harray[103][204], Harray[104][204], Harray[105][204], Harray[106][204], Harray[107][204], Harray[108][204], Harray[109][204], Harray[110][204], Harray[111][204], Harray[112][204], Harray[113][204], Harray[114][204], Harray[115][204], Harray[116][204], Harray[117][204], Harray[118][204], Harray[119][204], Harray[120][204], Harray[121][204], Harray[122][204], Harray[123][204], Harray[124][204], Harray[125][204], Harray[126][204], Harray[127][204]};
assign h_col_205 = {Harray[0][205], Harray[1][205], Harray[2][205], Harray[3][205], Harray[4][205], Harray[5][205], Harray[6][205], Harray[7][205], Harray[8][205], Harray[9][205], Harray[10][205], Harray[11][205], Harray[12][205], Harray[13][205], Harray[14][205], Harray[15][205], Harray[16][205], Harray[17][205], Harray[18][205], Harray[19][205], Harray[20][205], Harray[21][205], Harray[22][205], Harray[23][205], Harray[24][205], Harray[25][205], Harray[26][205], Harray[27][205], Harray[28][205], Harray[29][205], Harray[30][205], Harray[31][205], Harray[32][205], Harray[33][205], Harray[34][205], Harray[35][205], Harray[36][205], Harray[37][205], Harray[38][205], Harray[39][205], Harray[40][205], Harray[41][205], Harray[42][205], Harray[43][205], Harray[44][205], Harray[45][205], Harray[46][205], Harray[47][205], Harray[48][205], Harray[49][205], Harray[50][205], Harray[51][205], Harray[52][205], Harray[53][205], Harray[54][205], Harray[55][205], Harray[56][205], Harray[57][205], Harray[58][205], Harray[59][205], Harray[60][205], Harray[61][205], Harray[62][205], Harray[63][205], Harray[64][205], Harray[65][205], Harray[66][205], Harray[67][205], Harray[68][205], Harray[69][205], Harray[70][205], Harray[71][205], Harray[72][205], Harray[73][205], Harray[74][205], Harray[75][205], Harray[76][205], Harray[77][205], Harray[78][205], Harray[79][205], Harray[80][205], Harray[81][205], Harray[82][205], Harray[83][205], Harray[84][205], Harray[85][205], Harray[86][205], Harray[87][205], Harray[88][205], Harray[89][205], Harray[90][205], Harray[91][205], Harray[92][205], Harray[93][205], Harray[94][205], Harray[95][205], Harray[96][205], Harray[97][205], Harray[98][205], Harray[99][205], Harray[100][205], Harray[101][205], Harray[102][205], Harray[103][205], Harray[104][205], Harray[105][205], Harray[106][205], Harray[107][205], Harray[108][205], Harray[109][205], Harray[110][205], Harray[111][205], Harray[112][205], Harray[113][205], Harray[114][205], Harray[115][205], Harray[116][205], Harray[117][205], Harray[118][205], Harray[119][205], Harray[120][205], Harray[121][205], Harray[122][205], Harray[123][205], Harray[124][205], Harray[125][205], Harray[126][205], Harray[127][205]};
assign h_col_206 = {Harray[0][206], Harray[1][206], Harray[2][206], Harray[3][206], Harray[4][206], Harray[5][206], Harray[6][206], Harray[7][206], Harray[8][206], Harray[9][206], Harray[10][206], Harray[11][206], Harray[12][206], Harray[13][206], Harray[14][206], Harray[15][206], Harray[16][206], Harray[17][206], Harray[18][206], Harray[19][206], Harray[20][206], Harray[21][206], Harray[22][206], Harray[23][206], Harray[24][206], Harray[25][206], Harray[26][206], Harray[27][206], Harray[28][206], Harray[29][206], Harray[30][206], Harray[31][206], Harray[32][206], Harray[33][206], Harray[34][206], Harray[35][206], Harray[36][206], Harray[37][206], Harray[38][206], Harray[39][206], Harray[40][206], Harray[41][206], Harray[42][206], Harray[43][206], Harray[44][206], Harray[45][206], Harray[46][206], Harray[47][206], Harray[48][206], Harray[49][206], Harray[50][206], Harray[51][206], Harray[52][206], Harray[53][206], Harray[54][206], Harray[55][206], Harray[56][206], Harray[57][206], Harray[58][206], Harray[59][206], Harray[60][206], Harray[61][206], Harray[62][206], Harray[63][206], Harray[64][206], Harray[65][206], Harray[66][206], Harray[67][206], Harray[68][206], Harray[69][206], Harray[70][206], Harray[71][206], Harray[72][206], Harray[73][206], Harray[74][206], Harray[75][206], Harray[76][206], Harray[77][206], Harray[78][206], Harray[79][206], Harray[80][206], Harray[81][206], Harray[82][206], Harray[83][206], Harray[84][206], Harray[85][206], Harray[86][206], Harray[87][206], Harray[88][206], Harray[89][206], Harray[90][206], Harray[91][206], Harray[92][206], Harray[93][206], Harray[94][206], Harray[95][206], Harray[96][206], Harray[97][206], Harray[98][206], Harray[99][206], Harray[100][206], Harray[101][206], Harray[102][206], Harray[103][206], Harray[104][206], Harray[105][206], Harray[106][206], Harray[107][206], Harray[108][206], Harray[109][206], Harray[110][206], Harray[111][206], Harray[112][206], Harray[113][206], Harray[114][206], Harray[115][206], Harray[116][206], Harray[117][206], Harray[118][206], Harray[119][206], Harray[120][206], Harray[121][206], Harray[122][206], Harray[123][206], Harray[124][206], Harray[125][206], Harray[126][206], Harray[127][206]};
assign h_col_207 = {Harray[0][207], Harray[1][207], Harray[2][207], Harray[3][207], Harray[4][207], Harray[5][207], Harray[6][207], Harray[7][207], Harray[8][207], Harray[9][207], Harray[10][207], Harray[11][207], Harray[12][207], Harray[13][207], Harray[14][207], Harray[15][207], Harray[16][207], Harray[17][207], Harray[18][207], Harray[19][207], Harray[20][207], Harray[21][207], Harray[22][207], Harray[23][207], Harray[24][207], Harray[25][207], Harray[26][207], Harray[27][207], Harray[28][207], Harray[29][207], Harray[30][207], Harray[31][207], Harray[32][207], Harray[33][207], Harray[34][207], Harray[35][207], Harray[36][207], Harray[37][207], Harray[38][207], Harray[39][207], Harray[40][207], Harray[41][207], Harray[42][207], Harray[43][207], Harray[44][207], Harray[45][207], Harray[46][207], Harray[47][207], Harray[48][207], Harray[49][207], Harray[50][207], Harray[51][207], Harray[52][207], Harray[53][207], Harray[54][207], Harray[55][207], Harray[56][207], Harray[57][207], Harray[58][207], Harray[59][207], Harray[60][207], Harray[61][207], Harray[62][207], Harray[63][207], Harray[64][207], Harray[65][207], Harray[66][207], Harray[67][207], Harray[68][207], Harray[69][207], Harray[70][207], Harray[71][207], Harray[72][207], Harray[73][207], Harray[74][207], Harray[75][207], Harray[76][207], Harray[77][207], Harray[78][207], Harray[79][207], Harray[80][207], Harray[81][207], Harray[82][207], Harray[83][207], Harray[84][207], Harray[85][207], Harray[86][207], Harray[87][207], Harray[88][207], Harray[89][207], Harray[90][207], Harray[91][207], Harray[92][207], Harray[93][207], Harray[94][207], Harray[95][207], Harray[96][207], Harray[97][207], Harray[98][207], Harray[99][207], Harray[100][207], Harray[101][207], Harray[102][207], Harray[103][207], Harray[104][207], Harray[105][207], Harray[106][207], Harray[107][207], Harray[108][207], Harray[109][207], Harray[110][207], Harray[111][207], Harray[112][207], Harray[113][207], Harray[114][207], Harray[115][207], Harray[116][207], Harray[117][207], Harray[118][207], Harray[119][207], Harray[120][207], Harray[121][207], Harray[122][207], Harray[123][207], Harray[124][207], Harray[125][207], Harray[126][207], Harray[127][207]};
assign h_col_208 = {Harray[0][208], Harray[1][208], Harray[2][208], Harray[3][208], Harray[4][208], Harray[5][208], Harray[6][208], Harray[7][208], Harray[8][208], Harray[9][208], Harray[10][208], Harray[11][208], Harray[12][208], Harray[13][208], Harray[14][208], Harray[15][208], Harray[16][208], Harray[17][208], Harray[18][208], Harray[19][208], Harray[20][208], Harray[21][208], Harray[22][208], Harray[23][208], Harray[24][208], Harray[25][208], Harray[26][208], Harray[27][208], Harray[28][208], Harray[29][208], Harray[30][208], Harray[31][208], Harray[32][208], Harray[33][208], Harray[34][208], Harray[35][208], Harray[36][208], Harray[37][208], Harray[38][208], Harray[39][208], Harray[40][208], Harray[41][208], Harray[42][208], Harray[43][208], Harray[44][208], Harray[45][208], Harray[46][208], Harray[47][208], Harray[48][208], Harray[49][208], Harray[50][208], Harray[51][208], Harray[52][208], Harray[53][208], Harray[54][208], Harray[55][208], Harray[56][208], Harray[57][208], Harray[58][208], Harray[59][208], Harray[60][208], Harray[61][208], Harray[62][208], Harray[63][208], Harray[64][208], Harray[65][208], Harray[66][208], Harray[67][208], Harray[68][208], Harray[69][208], Harray[70][208], Harray[71][208], Harray[72][208], Harray[73][208], Harray[74][208], Harray[75][208], Harray[76][208], Harray[77][208], Harray[78][208], Harray[79][208], Harray[80][208], Harray[81][208], Harray[82][208], Harray[83][208], Harray[84][208], Harray[85][208], Harray[86][208], Harray[87][208], Harray[88][208], Harray[89][208], Harray[90][208], Harray[91][208], Harray[92][208], Harray[93][208], Harray[94][208], Harray[95][208], Harray[96][208], Harray[97][208], Harray[98][208], Harray[99][208], Harray[100][208], Harray[101][208], Harray[102][208], Harray[103][208], Harray[104][208], Harray[105][208], Harray[106][208], Harray[107][208], Harray[108][208], Harray[109][208], Harray[110][208], Harray[111][208], Harray[112][208], Harray[113][208], Harray[114][208], Harray[115][208], Harray[116][208], Harray[117][208], Harray[118][208], Harray[119][208], Harray[120][208], Harray[121][208], Harray[122][208], Harray[123][208], Harray[124][208], Harray[125][208], Harray[126][208], Harray[127][208]};
assign h_col_209 = {Harray[0][209], Harray[1][209], Harray[2][209], Harray[3][209], Harray[4][209], Harray[5][209], Harray[6][209], Harray[7][209], Harray[8][209], Harray[9][209], Harray[10][209], Harray[11][209], Harray[12][209], Harray[13][209], Harray[14][209], Harray[15][209], Harray[16][209], Harray[17][209], Harray[18][209], Harray[19][209], Harray[20][209], Harray[21][209], Harray[22][209], Harray[23][209], Harray[24][209], Harray[25][209], Harray[26][209], Harray[27][209], Harray[28][209], Harray[29][209], Harray[30][209], Harray[31][209], Harray[32][209], Harray[33][209], Harray[34][209], Harray[35][209], Harray[36][209], Harray[37][209], Harray[38][209], Harray[39][209], Harray[40][209], Harray[41][209], Harray[42][209], Harray[43][209], Harray[44][209], Harray[45][209], Harray[46][209], Harray[47][209], Harray[48][209], Harray[49][209], Harray[50][209], Harray[51][209], Harray[52][209], Harray[53][209], Harray[54][209], Harray[55][209], Harray[56][209], Harray[57][209], Harray[58][209], Harray[59][209], Harray[60][209], Harray[61][209], Harray[62][209], Harray[63][209], Harray[64][209], Harray[65][209], Harray[66][209], Harray[67][209], Harray[68][209], Harray[69][209], Harray[70][209], Harray[71][209], Harray[72][209], Harray[73][209], Harray[74][209], Harray[75][209], Harray[76][209], Harray[77][209], Harray[78][209], Harray[79][209], Harray[80][209], Harray[81][209], Harray[82][209], Harray[83][209], Harray[84][209], Harray[85][209], Harray[86][209], Harray[87][209], Harray[88][209], Harray[89][209], Harray[90][209], Harray[91][209], Harray[92][209], Harray[93][209], Harray[94][209], Harray[95][209], Harray[96][209], Harray[97][209], Harray[98][209], Harray[99][209], Harray[100][209], Harray[101][209], Harray[102][209], Harray[103][209], Harray[104][209], Harray[105][209], Harray[106][209], Harray[107][209], Harray[108][209], Harray[109][209], Harray[110][209], Harray[111][209], Harray[112][209], Harray[113][209], Harray[114][209], Harray[115][209], Harray[116][209], Harray[117][209], Harray[118][209], Harray[119][209], Harray[120][209], Harray[121][209], Harray[122][209], Harray[123][209], Harray[124][209], Harray[125][209], Harray[126][209], Harray[127][209]};
assign h_col_210 = {Harray[0][210], Harray[1][210], Harray[2][210], Harray[3][210], Harray[4][210], Harray[5][210], Harray[6][210], Harray[7][210], Harray[8][210], Harray[9][210], Harray[10][210], Harray[11][210], Harray[12][210], Harray[13][210], Harray[14][210], Harray[15][210], Harray[16][210], Harray[17][210], Harray[18][210], Harray[19][210], Harray[20][210], Harray[21][210], Harray[22][210], Harray[23][210], Harray[24][210], Harray[25][210], Harray[26][210], Harray[27][210], Harray[28][210], Harray[29][210], Harray[30][210], Harray[31][210], Harray[32][210], Harray[33][210], Harray[34][210], Harray[35][210], Harray[36][210], Harray[37][210], Harray[38][210], Harray[39][210], Harray[40][210], Harray[41][210], Harray[42][210], Harray[43][210], Harray[44][210], Harray[45][210], Harray[46][210], Harray[47][210], Harray[48][210], Harray[49][210], Harray[50][210], Harray[51][210], Harray[52][210], Harray[53][210], Harray[54][210], Harray[55][210], Harray[56][210], Harray[57][210], Harray[58][210], Harray[59][210], Harray[60][210], Harray[61][210], Harray[62][210], Harray[63][210], Harray[64][210], Harray[65][210], Harray[66][210], Harray[67][210], Harray[68][210], Harray[69][210], Harray[70][210], Harray[71][210], Harray[72][210], Harray[73][210], Harray[74][210], Harray[75][210], Harray[76][210], Harray[77][210], Harray[78][210], Harray[79][210], Harray[80][210], Harray[81][210], Harray[82][210], Harray[83][210], Harray[84][210], Harray[85][210], Harray[86][210], Harray[87][210], Harray[88][210], Harray[89][210], Harray[90][210], Harray[91][210], Harray[92][210], Harray[93][210], Harray[94][210], Harray[95][210], Harray[96][210], Harray[97][210], Harray[98][210], Harray[99][210], Harray[100][210], Harray[101][210], Harray[102][210], Harray[103][210], Harray[104][210], Harray[105][210], Harray[106][210], Harray[107][210], Harray[108][210], Harray[109][210], Harray[110][210], Harray[111][210], Harray[112][210], Harray[113][210], Harray[114][210], Harray[115][210], Harray[116][210], Harray[117][210], Harray[118][210], Harray[119][210], Harray[120][210], Harray[121][210], Harray[122][210], Harray[123][210], Harray[124][210], Harray[125][210], Harray[126][210], Harray[127][210]};
assign h_col_211 = {Harray[0][211], Harray[1][211], Harray[2][211], Harray[3][211], Harray[4][211], Harray[5][211], Harray[6][211], Harray[7][211], Harray[8][211], Harray[9][211], Harray[10][211], Harray[11][211], Harray[12][211], Harray[13][211], Harray[14][211], Harray[15][211], Harray[16][211], Harray[17][211], Harray[18][211], Harray[19][211], Harray[20][211], Harray[21][211], Harray[22][211], Harray[23][211], Harray[24][211], Harray[25][211], Harray[26][211], Harray[27][211], Harray[28][211], Harray[29][211], Harray[30][211], Harray[31][211], Harray[32][211], Harray[33][211], Harray[34][211], Harray[35][211], Harray[36][211], Harray[37][211], Harray[38][211], Harray[39][211], Harray[40][211], Harray[41][211], Harray[42][211], Harray[43][211], Harray[44][211], Harray[45][211], Harray[46][211], Harray[47][211], Harray[48][211], Harray[49][211], Harray[50][211], Harray[51][211], Harray[52][211], Harray[53][211], Harray[54][211], Harray[55][211], Harray[56][211], Harray[57][211], Harray[58][211], Harray[59][211], Harray[60][211], Harray[61][211], Harray[62][211], Harray[63][211], Harray[64][211], Harray[65][211], Harray[66][211], Harray[67][211], Harray[68][211], Harray[69][211], Harray[70][211], Harray[71][211], Harray[72][211], Harray[73][211], Harray[74][211], Harray[75][211], Harray[76][211], Harray[77][211], Harray[78][211], Harray[79][211], Harray[80][211], Harray[81][211], Harray[82][211], Harray[83][211], Harray[84][211], Harray[85][211], Harray[86][211], Harray[87][211], Harray[88][211], Harray[89][211], Harray[90][211], Harray[91][211], Harray[92][211], Harray[93][211], Harray[94][211], Harray[95][211], Harray[96][211], Harray[97][211], Harray[98][211], Harray[99][211], Harray[100][211], Harray[101][211], Harray[102][211], Harray[103][211], Harray[104][211], Harray[105][211], Harray[106][211], Harray[107][211], Harray[108][211], Harray[109][211], Harray[110][211], Harray[111][211], Harray[112][211], Harray[113][211], Harray[114][211], Harray[115][211], Harray[116][211], Harray[117][211], Harray[118][211], Harray[119][211], Harray[120][211], Harray[121][211], Harray[122][211], Harray[123][211], Harray[124][211], Harray[125][211], Harray[126][211], Harray[127][211]};
assign h_col_212 = {Harray[0][212], Harray[1][212], Harray[2][212], Harray[3][212], Harray[4][212], Harray[5][212], Harray[6][212], Harray[7][212], Harray[8][212], Harray[9][212], Harray[10][212], Harray[11][212], Harray[12][212], Harray[13][212], Harray[14][212], Harray[15][212], Harray[16][212], Harray[17][212], Harray[18][212], Harray[19][212], Harray[20][212], Harray[21][212], Harray[22][212], Harray[23][212], Harray[24][212], Harray[25][212], Harray[26][212], Harray[27][212], Harray[28][212], Harray[29][212], Harray[30][212], Harray[31][212], Harray[32][212], Harray[33][212], Harray[34][212], Harray[35][212], Harray[36][212], Harray[37][212], Harray[38][212], Harray[39][212], Harray[40][212], Harray[41][212], Harray[42][212], Harray[43][212], Harray[44][212], Harray[45][212], Harray[46][212], Harray[47][212], Harray[48][212], Harray[49][212], Harray[50][212], Harray[51][212], Harray[52][212], Harray[53][212], Harray[54][212], Harray[55][212], Harray[56][212], Harray[57][212], Harray[58][212], Harray[59][212], Harray[60][212], Harray[61][212], Harray[62][212], Harray[63][212], Harray[64][212], Harray[65][212], Harray[66][212], Harray[67][212], Harray[68][212], Harray[69][212], Harray[70][212], Harray[71][212], Harray[72][212], Harray[73][212], Harray[74][212], Harray[75][212], Harray[76][212], Harray[77][212], Harray[78][212], Harray[79][212], Harray[80][212], Harray[81][212], Harray[82][212], Harray[83][212], Harray[84][212], Harray[85][212], Harray[86][212], Harray[87][212], Harray[88][212], Harray[89][212], Harray[90][212], Harray[91][212], Harray[92][212], Harray[93][212], Harray[94][212], Harray[95][212], Harray[96][212], Harray[97][212], Harray[98][212], Harray[99][212], Harray[100][212], Harray[101][212], Harray[102][212], Harray[103][212], Harray[104][212], Harray[105][212], Harray[106][212], Harray[107][212], Harray[108][212], Harray[109][212], Harray[110][212], Harray[111][212], Harray[112][212], Harray[113][212], Harray[114][212], Harray[115][212], Harray[116][212], Harray[117][212], Harray[118][212], Harray[119][212], Harray[120][212], Harray[121][212], Harray[122][212], Harray[123][212], Harray[124][212], Harray[125][212], Harray[126][212], Harray[127][212]};
assign h_col_213 = {Harray[0][213], Harray[1][213], Harray[2][213], Harray[3][213], Harray[4][213], Harray[5][213], Harray[6][213], Harray[7][213], Harray[8][213], Harray[9][213], Harray[10][213], Harray[11][213], Harray[12][213], Harray[13][213], Harray[14][213], Harray[15][213], Harray[16][213], Harray[17][213], Harray[18][213], Harray[19][213], Harray[20][213], Harray[21][213], Harray[22][213], Harray[23][213], Harray[24][213], Harray[25][213], Harray[26][213], Harray[27][213], Harray[28][213], Harray[29][213], Harray[30][213], Harray[31][213], Harray[32][213], Harray[33][213], Harray[34][213], Harray[35][213], Harray[36][213], Harray[37][213], Harray[38][213], Harray[39][213], Harray[40][213], Harray[41][213], Harray[42][213], Harray[43][213], Harray[44][213], Harray[45][213], Harray[46][213], Harray[47][213], Harray[48][213], Harray[49][213], Harray[50][213], Harray[51][213], Harray[52][213], Harray[53][213], Harray[54][213], Harray[55][213], Harray[56][213], Harray[57][213], Harray[58][213], Harray[59][213], Harray[60][213], Harray[61][213], Harray[62][213], Harray[63][213], Harray[64][213], Harray[65][213], Harray[66][213], Harray[67][213], Harray[68][213], Harray[69][213], Harray[70][213], Harray[71][213], Harray[72][213], Harray[73][213], Harray[74][213], Harray[75][213], Harray[76][213], Harray[77][213], Harray[78][213], Harray[79][213], Harray[80][213], Harray[81][213], Harray[82][213], Harray[83][213], Harray[84][213], Harray[85][213], Harray[86][213], Harray[87][213], Harray[88][213], Harray[89][213], Harray[90][213], Harray[91][213], Harray[92][213], Harray[93][213], Harray[94][213], Harray[95][213], Harray[96][213], Harray[97][213], Harray[98][213], Harray[99][213], Harray[100][213], Harray[101][213], Harray[102][213], Harray[103][213], Harray[104][213], Harray[105][213], Harray[106][213], Harray[107][213], Harray[108][213], Harray[109][213], Harray[110][213], Harray[111][213], Harray[112][213], Harray[113][213], Harray[114][213], Harray[115][213], Harray[116][213], Harray[117][213], Harray[118][213], Harray[119][213], Harray[120][213], Harray[121][213], Harray[122][213], Harray[123][213], Harray[124][213], Harray[125][213], Harray[126][213], Harray[127][213]};
assign h_col_214 = {Harray[0][214], Harray[1][214], Harray[2][214], Harray[3][214], Harray[4][214], Harray[5][214], Harray[6][214], Harray[7][214], Harray[8][214], Harray[9][214], Harray[10][214], Harray[11][214], Harray[12][214], Harray[13][214], Harray[14][214], Harray[15][214], Harray[16][214], Harray[17][214], Harray[18][214], Harray[19][214], Harray[20][214], Harray[21][214], Harray[22][214], Harray[23][214], Harray[24][214], Harray[25][214], Harray[26][214], Harray[27][214], Harray[28][214], Harray[29][214], Harray[30][214], Harray[31][214], Harray[32][214], Harray[33][214], Harray[34][214], Harray[35][214], Harray[36][214], Harray[37][214], Harray[38][214], Harray[39][214], Harray[40][214], Harray[41][214], Harray[42][214], Harray[43][214], Harray[44][214], Harray[45][214], Harray[46][214], Harray[47][214], Harray[48][214], Harray[49][214], Harray[50][214], Harray[51][214], Harray[52][214], Harray[53][214], Harray[54][214], Harray[55][214], Harray[56][214], Harray[57][214], Harray[58][214], Harray[59][214], Harray[60][214], Harray[61][214], Harray[62][214], Harray[63][214], Harray[64][214], Harray[65][214], Harray[66][214], Harray[67][214], Harray[68][214], Harray[69][214], Harray[70][214], Harray[71][214], Harray[72][214], Harray[73][214], Harray[74][214], Harray[75][214], Harray[76][214], Harray[77][214], Harray[78][214], Harray[79][214], Harray[80][214], Harray[81][214], Harray[82][214], Harray[83][214], Harray[84][214], Harray[85][214], Harray[86][214], Harray[87][214], Harray[88][214], Harray[89][214], Harray[90][214], Harray[91][214], Harray[92][214], Harray[93][214], Harray[94][214], Harray[95][214], Harray[96][214], Harray[97][214], Harray[98][214], Harray[99][214], Harray[100][214], Harray[101][214], Harray[102][214], Harray[103][214], Harray[104][214], Harray[105][214], Harray[106][214], Harray[107][214], Harray[108][214], Harray[109][214], Harray[110][214], Harray[111][214], Harray[112][214], Harray[113][214], Harray[114][214], Harray[115][214], Harray[116][214], Harray[117][214], Harray[118][214], Harray[119][214], Harray[120][214], Harray[121][214], Harray[122][214], Harray[123][214], Harray[124][214], Harray[125][214], Harray[126][214], Harray[127][214]};
assign h_col_215 = {Harray[0][215], Harray[1][215], Harray[2][215], Harray[3][215], Harray[4][215], Harray[5][215], Harray[6][215], Harray[7][215], Harray[8][215], Harray[9][215], Harray[10][215], Harray[11][215], Harray[12][215], Harray[13][215], Harray[14][215], Harray[15][215], Harray[16][215], Harray[17][215], Harray[18][215], Harray[19][215], Harray[20][215], Harray[21][215], Harray[22][215], Harray[23][215], Harray[24][215], Harray[25][215], Harray[26][215], Harray[27][215], Harray[28][215], Harray[29][215], Harray[30][215], Harray[31][215], Harray[32][215], Harray[33][215], Harray[34][215], Harray[35][215], Harray[36][215], Harray[37][215], Harray[38][215], Harray[39][215], Harray[40][215], Harray[41][215], Harray[42][215], Harray[43][215], Harray[44][215], Harray[45][215], Harray[46][215], Harray[47][215], Harray[48][215], Harray[49][215], Harray[50][215], Harray[51][215], Harray[52][215], Harray[53][215], Harray[54][215], Harray[55][215], Harray[56][215], Harray[57][215], Harray[58][215], Harray[59][215], Harray[60][215], Harray[61][215], Harray[62][215], Harray[63][215], Harray[64][215], Harray[65][215], Harray[66][215], Harray[67][215], Harray[68][215], Harray[69][215], Harray[70][215], Harray[71][215], Harray[72][215], Harray[73][215], Harray[74][215], Harray[75][215], Harray[76][215], Harray[77][215], Harray[78][215], Harray[79][215], Harray[80][215], Harray[81][215], Harray[82][215], Harray[83][215], Harray[84][215], Harray[85][215], Harray[86][215], Harray[87][215], Harray[88][215], Harray[89][215], Harray[90][215], Harray[91][215], Harray[92][215], Harray[93][215], Harray[94][215], Harray[95][215], Harray[96][215], Harray[97][215], Harray[98][215], Harray[99][215], Harray[100][215], Harray[101][215], Harray[102][215], Harray[103][215], Harray[104][215], Harray[105][215], Harray[106][215], Harray[107][215], Harray[108][215], Harray[109][215], Harray[110][215], Harray[111][215], Harray[112][215], Harray[113][215], Harray[114][215], Harray[115][215], Harray[116][215], Harray[117][215], Harray[118][215], Harray[119][215], Harray[120][215], Harray[121][215], Harray[122][215], Harray[123][215], Harray[124][215], Harray[125][215], Harray[126][215], Harray[127][215]};
assign h_col_216 = {Harray[0][216], Harray[1][216], Harray[2][216], Harray[3][216], Harray[4][216], Harray[5][216], Harray[6][216], Harray[7][216], Harray[8][216], Harray[9][216], Harray[10][216], Harray[11][216], Harray[12][216], Harray[13][216], Harray[14][216], Harray[15][216], Harray[16][216], Harray[17][216], Harray[18][216], Harray[19][216], Harray[20][216], Harray[21][216], Harray[22][216], Harray[23][216], Harray[24][216], Harray[25][216], Harray[26][216], Harray[27][216], Harray[28][216], Harray[29][216], Harray[30][216], Harray[31][216], Harray[32][216], Harray[33][216], Harray[34][216], Harray[35][216], Harray[36][216], Harray[37][216], Harray[38][216], Harray[39][216], Harray[40][216], Harray[41][216], Harray[42][216], Harray[43][216], Harray[44][216], Harray[45][216], Harray[46][216], Harray[47][216], Harray[48][216], Harray[49][216], Harray[50][216], Harray[51][216], Harray[52][216], Harray[53][216], Harray[54][216], Harray[55][216], Harray[56][216], Harray[57][216], Harray[58][216], Harray[59][216], Harray[60][216], Harray[61][216], Harray[62][216], Harray[63][216], Harray[64][216], Harray[65][216], Harray[66][216], Harray[67][216], Harray[68][216], Harray[69][216], Harray[70][216], Harray[71][216], Harray[72][216], Harray[73][216], Harray[74][216], Harray[75][216], Harray[76][216], Harray[77][216], Harray[78][216], Harray[79][216], Harray[80][216], Harray[81][216], Harray[82][216], Harray[83][216], Harray[84][216], Harray[85][216], Harray[86][216], Harray[87][216], Harray[88][216], Harray[89][216], Harray[90][216], Harray[91][216], Harray[92][216], Harray[93][216], Harray[94][216], Harray[95][216], Harray[96][216], Harray[97][216], Harray[98][216], Harray[99][216], Harray[100][216], Harray[101][216], Harray[102][216], Harray[103][216], Harray[104][216], Harray[105][216], Harray[106][216], Harray[107][216], Harray[108][216], Harray[109][216], Harray[110][216], Harray[111][216], Harray[112][216], Harray[113][216], Harray[114][216], Harray[115][216], Harray[116][216], Harray[117][216], Harray[118][216], Harray[119][216], Harray[120][216], Harray[121][216], Harray[122][216], Harray[123][216], Harray[124][216], Harray[125][216], Harray[126][216], Harray[127][216]};
assign h_col_217 = {Harray[0][217], Harray[1][217], Harray[2][217], Harray[3][217], Harray[4][217], Harray[5][217], Harray[6][217], Harray[7][217], Harray[8][217], Harray[9][217], Harray[10][217], Harray[11][217], Harray[12][217], Harray[13][217], Harray[14][217], Harray[15][217], Harray[16][217], Harray[17][217], Harray[18][217], Harray[19][217], Harray[20][217], Harray[21][217], Harray[22][217], Harray[23][217], Harray[24][217], Harray[25][217], Harray[26][217], Harray[27][217], Harray[28][217], Harray[29][217], Harray[30][217], Harray[31][217], Harray[32][217], Harray[33][217], Harray[34][217], Harray[35][217], Harray[36][217], Harray[37][217], Harray[38][217], Harray[39][217], Harray[40][217], Harray[41][217], Harray[42][217], Harray[43][217], Harray[44][217], Harray[45][217], Harray[46][217], Harray[47][217], Harray[48][217], Harray[49][217], Harray[50][217], Harray[51][217], Harray[52][217], Harray[53][217], Harray[54][217], Harray[55][217], Harray[56][217], Harray[57][217], Harray[58][217], Harray[59][217], Harray[60][217], Harray[61][217], Harray[62][217], Harray[63][217], Harray[64][217], Harray[65][217], Harray[66][217], Harray[67][217], Harray[68][217], Harray[69][217], Harray[70][217], Harray[71][217], Harray[72][217], Harray[73][217], Harray[74][217], Harray[75][217], Harray[76][217], Harray[77][217], Harray[78][217], Harray[79][217], Harray[80][217], Harray[81][217], Harray[82][217], Harray[83][217], Harray[84][217], Harray[85][217], Harray[86][217], Harray[87][217], Harray[88][217], Harray[89][217], Harray[90][217], Harray[91][217], Harray[92][217], Harray[93][217], Harray[94][217], Harray[95][217], Harray[96][217], Harray[97][217], Harray[98][217], Harray[99][217], Harray[100][217], Harray[101][217], Harray[102][217], Harray[103][217], Harray[104][217], Harray[105][217], Harray[106][217], Harray[107][217], Harray[108][217], Harray[109][217], Harray[110][217], Harray[111][217], Harray[112][217], Harray[113][217], Harray[114][217], Harray[115][217], Harray[116][217], Harray[117][217], Harray[118][217], Harray[119][217], Harray[120][217], Harray[121][217], Harray[122][217], Harray[123][217], Harray[124][217], Harray[125][217], Harray[126][217], Harray[127][217]};
assign h_col_218 = {Harray[0][218], Harray[1][218], Harray[2][218], Harray[3][218], Harray[4][218], Harray[5][218], Harray[6][218], Harray[7][218], Harray[8][218], Harray[9][218], Harray[10][218], Harray[11][218], Harray[12][218], Harray[13][218], Harray[14][218], Harray[15][218], Harray[16][218], Harray[17][218], Harray[18][218], Harray[19][218], Harray[20][218], Harray[21][218], Harray[22][218], Harray[23][218], Harray[24][218], Harray[25][218], Harray[26][218], Harray[27][218], Harray[28][218], Harray[29][218], Harray[30][218], Harray[31][218], Harray[32][218], Harray[33][218], Harray[34][218], Harray[35][218], Harray[36][218], Harray[37][218], Harray[38][218], Harray[39][218], Harray[40][218], Harray[41][218], Harray[42][218], Harray[43][218], Harray[44][218], Harray[45][218], Harray[46][218], Harray[47][218], Harray[48][218], Harray[49][218], Harray[50][218], Harray[51][218], Harray[52][218], Harray[53][218], Harray[54][218], Harray[55][218], Harray[56][218], Harray[57][218], Harray[58][218], Harray[59][218], Harray[60][218], Harray[61][218], Harray[62][218], Harray[63][218], Harray[64][218], Harray[65][218], Harray[66][218], Harray[67][218], Harray[68][218], Harray[69][218], Harray[70][218], Harray[71][218], Harray[72][218], Harray[73][218], Harray[74][218], Harray[75][218], Harray[76][218], Harray[77][218], Harray[78][218], Harray[79][218], Harray[80][218], Harray[81][218], Harray[82][218], Harray[83][218], Harray[84][218], Harray[85][218], Harray[86][218], Harray[87][218], Harray[88][218], Harray[89][218], Harray[90][218], Harray[91][218], Harray[92][218], Harray[93][218], Harray[94][218], Harray[95][218], Harray[96][218], Harray[97][218], Harray[98][218], Harray[99][218], Harray[100][218], Harray[101][218], Harray[102][218], Harray[103][218], Harray[104][218], Harray[105][218], Harray[106][218], Harray[107][218], Harray[108][218], Harray[109][218], Harray[110][218], Harray[111][218], Harray[112][218], Harray[113][218], Harray[114][218], Harray[115][218], Harray[116][218], Harray[117][218], Harray[118][218], Harray[119][218], Harray[120][218], Harray[121][218], Harray[122][218], Harray[123][218], Harray[124][218], Harray[125][218], Harray[126][218], Harray[127][218]};
assign h_col_219 = {Harray[0][219], Harray[1][219], Harray[2][219], Harray[3][219], Harray[4][219], Harray[5][219], Harray[6][219], Harray[7][219], Harray[8][219], Harray[9][219], Harray[10][219], Harray[11][219], Harray[12][219], Harray[13][219], Harray[14][219], Harray[15][219], Harray[16][219], Harray[17][219], Harray[18][219], Harray[19][219], Harray[20][219], Harray[21][219], Harray[22][219], Harray[23][219], Harray[24][219], Harray[25][219], Harray[26][219], Harray[27][219], Harray[28][219], Harray[29][219], Harray[30][219], Harray[31][219], Harray[32][219], Harray[33][219], Harray[34][219], Harray[35][219], Harray[36][219], Harray[37][219], Harray[38][219], Harray[39][219], Harray[40][219], Harray[41][219], Harray[42][219], Harray[43][219], Harray[44][219], Harray[45][219], Harray[46][219], Harray[47][219], Harray[48][219], Harray[49][219], Harray[50][219], Harray[51][219], Harray[52][219], Harray[53][219], Harray[54][219], Harray[55][219], Harray[56][219], Harray[57][219], Harray[58][219], Harray[59][219], Harray[60][219], Harray[61][219], Harray[62][219], Harray[63][219], Harray[64][219], Harray[65][219], Harray[66][219], Harray[67][219], Harray[68][219], Harray[69][219], Harray[70][219], Harray[71][219], Harray[72][219], Harray[73][219], Harray[74][219], Harray[75][219], Harray[76][219], Harray[77][219], Harray[78][219], Harray[79][219], Harray[80][219], Harray[81][219], Harray[82][219], Harray[83][219], Harray[84][219], Harray[85][219], Harray[86][219], Harray[87][219], Harray[88][219], Harray[89][219], Harray[90][219], Harray[91][219], Harray[92][219], Harray[93][219], Harray[94][219], Harray[95][219], Harray[96][219], Harray[97][219], Harray[98][219], Harray[99][219], Harray[100][219], Harray[101][219], Harray[102][219], Harray[103][219], Harray[104][219], Harray[105][219], Harray[106][219], Harray[107][219], Harray[108][219], Harray[109][219], Harray[110][219], Harray[111][219], Harray[112][219], Harray[113][219], Harray[114][219], Harray[115][219], Harray[116][219], Harray[117][219], Harray[118][219], Harray[119][219], Harray[120][219], Harray[121][219], Harray[122][219], Harray[123][219], Harray[124][219], Harray[125][219], Harray[126][219], Harray[127][219]};
assign h_col_220 = {Harray[0][220], Harray[1][220], Harray[2][220], Harray[3][220], Harray[4][220], Harray[5][220], Harray[6][220], Harray[7][220], Harray[8][220], Harray[9][220], Harray[10][220], Harray[11][220], Harray[12][220], Harray[13][220], Harray[14][220], Harray[15][220], Harray[16][220], Harray[17][220], Harray[18][220], Harray[19][220], Harray[20][220], Harray[21][220], Harray[22][220], Harray[23][220], Harray[24][220], Harray[25][220], Harray[26][220], Harray[27][220], Harray[28][220], Harray[29][220], Harray[30][220], Harray[31][220], Harray[32][220], Harray[33][220], Harray[34][220], Harray[35][220], Harray[36][220], Harray[37][220], Harray[38][220], Harray[39][220], Harray[40][220], Harray[41][220], Harray[42][220], Harray[43][220], Harray[44][220], Harray[45][220], Harray[46][220], Harray[47][220], Harray[48][220], Harray[49][220], Harray[50][220], Harray[51][220], Harray[52][220], Harray[53][220], Harray[54][220], Harray[55][220], Harray[56][220], Harray[57][220], Harray[58][220], Harray[59][220], Harray[60][220], Harray[61][220], Harray[62][220], Harray[63][220], Harray[64][220], Harray[65][220], Harray[66][220], Harray[67][220], Harray[68][220], Harray[69][220], Harray[70][220], Harray[71][220], Harray[72][220], Harray[73][220], Harray[74][220], Harray[75][220], Harray[76][220], Harray[77][220], Harray[78][220], Harray[79][220], Harray[80][220], Harray[81][220], Harray[82][220], Harray[83][220], Harray[84][220], Harray[85][220], Harray[86][220], Harray[87][220], Harray[88][220], Harray[89][220], Harray[90][220], Harray[91][220], Harray[92][220], Harray[93][220], Harray[94][220], Harray[95][220], Harray[96][220], Harray[97][220], Harray[98][220], Harray[99][220], Harray[100][220], Harray[101][220], Harray[102][220], Harray[103][220], Harray[104][220], Harray[105][220], Harray[106][220], Harray[107][220], Harray[108][220], Harray[109][220], Harray[110][220], Harray[111][220], Harray[112][220], Harray[113][220], Harray[114][220], Harray[115][220], Harray[116][220], Harray[117][220], Harray[118][220], Harray[119][220], Harray[120][220], Harray[121][220], Harray[122][220], Harray[123][220], Harray[124][220], Harray[125][220], Harray[126][220], Harray[127][220]};
assign h_col_221 = {Harray[0][221], Harray[1][221], Harray[2][221], Harray[3][221], Harray[4][221], Harray[5][221], Harray[6][221], Harray[7][221], Harray[8][221], Harray[9][221], Harray[10][221], Harray[11][221], Harray[12][221], Harray[13][221], Harray[14][221], Harray[15][221], Harray[16][221], Harray[17][221], Harray[18][221], Harray[19][221], Harray[20][221], Harray[21][221], Harray[22][221], Harray[23][221], Harray[24][221], Harray[25][221], Harray[26][221], Harray[27][221], Harray[28][221], Harray[29][221], Harray[30][221], Harray[31][221], Harray[32][221], Harray[33][221], Harray[34][221], Harray[35][221], Harray[36][221], Harray[37][221], Harray[38][221], Harray[39][221], Harray[40][221], Harray[41][221], Harray[42][221], Harray[43][221], Harray[44][221], Harray[45][221], Harray[46][221], Harray[47][221], Harray[48][221], Harray[49][221], Harray[50][221], Harray[51][221], Harray[52][221], Harray[53][221], Harray[54][221], Harray[55][221], Harray[56][221], Harray[57][221], Harray[58][221], Harray[59][221], Harray[60][221], Harray[61][221], Harray[62][221], Harray[63][221], Harray[64][221], Harray[65][221], Harray[66][221], Harray[67][221], Harray[68][221], Harray[69][221], Harray[70][221], Harray[71][221], Harray[72][221], Harray[73][221], Harray[74][221], Harray[75][221], Harray[76][221], Harray[77][221], Harray[78][221], Harray[79][221], Harray[80][221], Harray[81][221], Harray[82][221], Harray[83][221], Harray[84][221], Harray[85][221], Harray[86][221], Harray[87][221], Harray[88][221], Harray[89][221], Harray[90][221], Harray[91][221], Harray[92][221], Harray[93][221], Harray[94][221], Harray[95][221], Harray[96][221], Harray[97][221], Harray[98][221], Harray[99][221], Harray[100][221], Harray[101][221], Harray[102][221], Harray[103][221], Harray[104][221], Harray[105][221], Harray[106][221], Harray[107][221], Harray[108][221], Harray[109][221], Harray[110][221], Harray[111][221], Harray[112][221], Harray[113][221], Harray[114][221], Harray[115][221], Harray[116][221], Harray[117][221], Harray[118][221], Harray[119][221], Harray[120][221], Harray[121][221], Harray[122][221], Harray[123][221], Harray[124][221], Harray[125][221], Harray[126][221], Harray[127][221]};
assign h_col_222 = {Harray[0][222], Harray[1][222], Harray[2][222], Harray[3][222], Harray[4][222], Harray[5][222], Harray[6][222], Harray[7][222], Harray[8][222], Harray[9][222], Harray[10][222], Harray[11][222], Harray[12][222], Harray[13][222], Harray[14][222], Harray[15][222], Harray[16][222], Harray[17][222], Harray[18][222], Harray[19][222], Harray[20][222], Harray[21][222], Harray[22][222], Harray[23][222], Harray[24][222], Harray[25][222], Harray[26][222], Harray[27][222], Harray[28][222], Harray[29][222], Harray[30][222], Harray[31][222], Harray[32][222], Harray[33][222], Harray[34][222], Harray[35][222], Harray[36][222], Harray[37][222], Harray[38][222], Harray[39][222], Harray[40][222], Harray[41][222], Harray[42][222], Harray[43][222], Harray[44][222], Harray[45][222], Harray[46][222], Harray[47][222], Harray[48][222], Harray[49][222], Harray[50][222], Harray[51][222], Harray[52][222], Harray[53][222], Harray[54][222], Harray[55][222], Harray[56][222], Harray[57][222], Harray[58][222], Harray[59][222], Harray[60][222], Harray[61][222], Harray[62][222], Harray[63][222], Harray[64][222], Harray[65][222], Harray[66][222], Harray[67][222], Harray[68][222], Harray[69][222], Harray[70][222], Harray[71][222], Harray[72][222], Harray[73][222], Harray[74][222], Harray[75][222], Harray[76][222], Harray[77][222], Harray[78][222], Harray[79][222], Harray[80][222], Harray[81][222], Harray[82][222], Harray[83][222], Harray[84][222], Harray[85][222], Harray[86][222], Harray[87][222], Harray[88][222], Harray[89][222], Harray[90][222], Harray[91][222], Harray[92][222], Harray[93][222], Harray[94][222], Harray[95][222], Harray[96][222], Harray[97][222], Harray[98][222], Harray[99][222], Harray[100][222], Harray[101][222], Harray[102][222], Harray[103][222], Harray[104][222], Harray[105][222], Harray[106][222], Harray[107][222], Harray[108][222], Harray[109][222], Harray[110][222], Harray[111][222], Harray[112][222], Harray[113][222], Harray[114][222], Harray[115][222], Harray[116][222], Harray[117][222], Harray[118][222], Harray[119][222], Harray[120][222], Harray[121][222], Harray[122][222], Harray[123][222], Harray[124][222], Harray[125][222], Harray[126][222], Harray[127][222]};
assign h_col_223 = {Harray[0][223], Harray[1][223], Harray[2][223], Harray[3][223], Harray[4][223], Harray[5][223], Harray[6][223], Harray[7][223], Harray[8][223], Harray[9][223], Harray[10][223], Harray[11][223], Harray[12][223], Harray[13][223], Harray[14][223], Harray[15][223], Harray[16][223], Harray[17][223], Harray[18][223], Harray[19][223], Harray[20][223], Harray[21][223], Harray[22][223], Harray[23][223], Harray[24][223], Harray[25][223], Harray[26][223], Harray[27][223], Harray[28][223], Harray[29][223], Harray[30][223], Harray[31][223], Harray[32][223], Harray[33][223], Harray[34][223], Harray[35][223], Harray[36][223], Harray[37][223], Harray[38][223], Harray[39][223], Harray[40][223], Harray[41][223], Harray[42][223], Harray[43][223], Harray[44][223], Harray[45][223], Harray[46][223], Harray[47][223], Harray[48][223], Harray[49][223], Harray[50][223], Harray[51][223], Harray[52][223], Harray[53][223], Harray[54][223], Harray[55][223], Harray[56][223], Harray[57][223], Harray[58][223], Harray[59][223], Harray[60][223], Harray[61][223], Harray[62][223], Harray[63][223], Harray[64][223], Harray[65][223], Harray[66][223], Harray[67][223], Harray[68][223], Harray[69][223], Harray[70][223], Harray[71][223], Harray[72][223], Harray[73][223], Harray[74][223], Harray[75][223], Harray[76][223], Harray[77][223], Harray[78][223], Harray[79][223], Harray[80][223], Harray[81][223], Harray[82][223], Harray[83][223], Harray[84][223], Harray[85][223], Harray[86][223], Harray[87][223], Harray[88][223], Harray[89][223], Harray[90][223], Harray[91][223], Harray[92][223], Harray[93][223], Harray[94][223], Harray[95][223], Harray[96][223], Harray[97][223], Harray[98][223], Harray[99][223], Harray[100][223], Harray[101][223], Harray[102][223], Harray[103][223], Harray[104][223], Harray[105][223], Harray[106][223], Harray[107][223], Harray[108][223], Harray[109][223], Harray[110][223], Harray[111][223], Harray[112][223], Harray[113][223], Harray[114][223], Harray[115][223], Harray[116][223], Harray[117][223], Harray[118][223], Harray[119][223], Harray[120][223], Harray[121][223], Harray[122][223], Harray[123][223], Harray[124][223], Harray[125][223], Harray[126][223], Harray[127][223]};
assign h_col_224 = {Harray[0][224], Harray[1][224], Harray[2][224], Harray[3][224], Harray[4][224], Harray[5][224], Harray[6][224], Harray[7][224], Harray[8][224], Harray[9][224], Harray[10][224], Harray[11][224], Harray[12][224], Harray[13][224], Harray[14][224], Harray[15][224], Harray[16][224], Harray[17][224], Harray[18][224], Harray[19][224], Harray[20][224], Harray[21][224], Harray[22][224], Harray[23][224], Harray[24][224], Harray[25][224], Harray[26][224], Harray[27][224], Harray[28][224], Harray[29][224], Harray[30][224], Harray[31][224], Harray[32][224], Harray[33][224], Harray[34][224], Harray[35][224], Harray[36][224], Harray[37][224], Harray[38][224], Harray[39][224], Harray[40][224], Harray[41][224], Harray[42][224], Harray[43][224], Harray[44][224], Harray[45][224], Harray[46][224], Harray[47][224], Harray[48][224], Harray[49][224], Harray[50][224], Harray[51][224], Harray[52][224], Harray[53][224], Harray[54][224], Harray[55][224], Harray[56][224], Harray[57][224], Harray[58][224], Harray[59][224], Harray[60][224], Harray[61][224], Harray[62][224], Harray[63][224], Harray[64][224], Harray[65][224], Harray[66][224], Harray[67][224], Harray[68][224], Harray[69][224], Harray[70][224], Harray[71][224], Harray[72][224], Harray[73][224], Harray[74][224], Harray[75][224], Harray[76][224], Harray[77][224], Harray[78][224], Harray[79][224], Harray[80][224], Harray[81][224], Harray[82][224], Harray[83][224], Harray[84][224], Harray[85][224], Harray[86][224], Harray[87][224], Harray[88][224], Harray[89][224], Harray[90][224], Harray[91][224], Harray[92][224], Harray[93][224], Harray[94][224], Harray[95][224], Harray[96][224], Harray[97][224], Harray[98][224], Harray[99][224], Harray[100][224], Harray[101][224], Harray[102][224], Harray[103][224], Harray[104][224], Harray[105][224], Harray[106][224], Harray[107][224], Harray[108][224], Harray[109][224], Harray[110][224], Harray[111][224], Harray[112][224], Harray[113][224], Harray[114][224], Harray[115][224], Harray[116][224], Harray[117][224], Harray[118][224], Harray[119][224], Harray[120][224], Harray[121][224], Harray[122][224], Harray[123][224], Harray[124][224], Harray[125][224], Harray[126][224], Harray[127][224]};
assign h_col_225 = {Harray[0][225], Harray[1][225], Harray[2][225], Harray[3][225], Harray[4][225], Harray[5][225], Harray[6][225], Harray[7][225], Harray[8][225], Harray[9][225], Harray[10][225], Harray[11][225], Harray[12][225], Harray[13][225], Harray[14][225], Harray[15][225], Harray[16][225], Harray[17][225], Harray[18][225], Harray[19][225], Harray[20][225], Harray[21][225], Harray[22][225], Harray[23][225], Harray[24][225], Harray[25][225], Harray[26][225], Harray[27][225], Harray[28][225], Harray[29][225], Harray[30][225], Harray[31][225], Harray[32][225], Harray[33][225], Harray[34][225], Harray[35][225], Harray[36][225], Harray[37][225], Harray[38][225], Harray[39][225], Harray[40][225], Harray[41][225], Harray[42][225], Harray[43][225], Harray[44][225], Harray[45][225], Harray[46][225], Harray[47][225], Harray[48][225], Harray[49][225], Harray[50][225], Harray[51][225], Harray[52][225], Harray[53][225], Harray[54][225], Harray[55][225], Harray[56][225], Harray[57][225], Harray[58][225], Harray[59][225], Harray[60][225], Harray[61][225], Harray[62][225], Harray[63][225], Harray[64][225], Harray[65][225], Harray[66][225], Harray[67][225], Harray[68][225], Harray[69][225], Harray[70][225], Harray[71][225], Harray[72][225], Harray[73][225], Harray[74][225], Harray[75][225], Harray[76][225], Harray[77][225], Harray[78][225], Harray[79][225], Harray[80][225], Harray[81][225], Harray[82][225], Harray[83][225], Harray[84][225], Harray[85][225], Harray[86][225], Harray[87][225], Harray[88][225], Harray[89][225], Harray[90][225], Harray[91][225], Harray[92][225], Harray[93][225], Harray[94][225], Harray[95][225], Harray[96][225], Harray[97][225], Harray[98][225], Harray[99][225], Harray[100][225], Harray[101][225], Harray[102][225], Harray[103][225], Harray[104][225], Harray[105][225], Harray[106][225], Harray[107][225], Harray[108][225], Harray[109][225], Harray[110][225], Harray[111][225], Harray[112][225], Harray[113][225], Harray[114][225], Harray[115][225], Harray[116][225], Harray[117][225], Harray[118][225], Harray[119][225], Harray[120][225], Harray[121][225], Harray[122][225], Harray[123][225], Harray[124][225], Harray[125][225], Harray[126][225], Harray[127][225]};
assign h_col_226 = {Harray[0][226], Harray[1][226], Harray[2][226], Harray[3][226], Harray[4][226], Harray[5][226], Harray[6][226], Harray[7][226], Harray[8][226], Harray[9][226], Harray[10][226], Harray[11][226], Harray[12][226], Harray[13][226], Harray[14][226], Harray[15][226], Harray[16][226], Harray[17][226], Harray[18][226], Harray[19][226], Harray[20][226], Harray[21][226], Harray[22][226], Harray[23][226], Harray[24][226], Harray[25][226], Harray[26][226], Harray[27][226], Harray[28][226], Harray[29][226], Harray[30][226], Harray[31][226], Harray[32][226], Harray[33][226], Harray[34][226], Harray[35][226], Harray[36][226], Harray[37][226], Harray[38][226], Harray[39][226], Harray[40][226], Harray[41][226], Harray[42][226], Harray[43][226], Harray[44][226], Harray[45][226], Harray[46][226], Harray[47][226], Harray[48][226], Harray[49][226], Harray[50][226], Harray[51][226], Harray[52][226], Harray[53][226], Harray[54][226], Harray[55][226], Harray[56][226], Harray[57][226], Harray[58][226], Harray[59][226], Harray[60][226], Harray[61][226], Harray[62][226], Harray[63][226], Harray[64][226], Harray[65][226], Harray[66][226], Harray[67][226], Harray[68][226], Harray[69][226], Harray[70][226], Harray[71][226], Harray[72][226], Harray[73][226], Harray[74][226], Harray[75][226], Harray[76][226], Harray[77][226], Harray[78][226], Harray[79][226], Harray[80][226], Harray[81][226], Harray[82][226], Harray[83][226], Harray[84][226], Harray[85][226], Harray[86][226], Harray[87][226], Harray[88][226], Harray[89][226], Harray[90][226], Harray[91][226], Harray[92][226], Harray[93][226], Harray[94][226], Harray[95][226], Harray[96][226], Harray[97][226], Harray[98][226], Harray[99][226], Harray[100][226], Harray[101][226], Harray[102][226], Harray[103][226], Harray[104][226], Harray[105][226], Harray[106][226], Harray[107][226], Harray[108][226], Harray[109][226], Harray[110][226], Harray[111][226], Harray[112][226], Harray[113][226], Harray[114][226], Harray[115][226], Harray[116][226], Harray[117][226], Harray[118][226], Harray[119][226], Harray[120][226], Harray[121][226], Harray[122][226], Harray[123][226], Harray[124][226], Harray[125][226], Harray[126][226], Harray[127][226]};
assign h_col_227 = {Harray[0][227], Harray[1][227], Harray[2][227], Harray[3][227], Harray[4][227], Harray[5][227], Harray[6][227], Harray[7][227], Harray[8][227], Harray[9][227], Harray[10][227], Harray[11][227], Harray[12][227], Harray[13][227], Harray[14][227], Harray[15][227], Harray[16][227], Harray[17][227], Harray[18][227], Harray[19][227], Harray[20][227], Harray[21][227], Harray[22][227], Harray[23][227], Harray[24][227], Harray[25][227], Harray[26][227], Harray[27][227], Harray[28][227], Harray[29][227], Harray[30][227], Harray[31][227], Harray[32][227], Harray[33][227], Harray[34][227], Harray[35][227], Harray[36][227], Harray[37][227], Harray[38][227], Harray[39][227], Harray[40][227], Harray[41][227], Harray[42][227], Harray[43][227], Harray[44][227], Harray[45][227], Harray[46][227], Harray[47][227], Harray[48][227], Harray[49][227], Harray[50][227], Harray[51][227], Harray[52][227], Harray[53][227], Harray[54][227], Harray[55][227], Harray[56][227], Harray[57][227], Harray[58][227], Harray[59][227], Harray[60][227], Harray[61][227], Harray[62][227], Harray[63][227], Harray[64][227], Harray[65][227], Harray[66][227], Harray[67][227], Harray[68][227], Harray[69][227], Harray[70][227], Harray[71][227], Harray[72][227], Harray[73][227], Harray[74][227], Harray[75][227], Harray[76][227], Harray[77][227], Harray[78][227], Harray[79][227], Harray[80][227], Harray[81][227], Harray[82][227], Harray[83][227], Harray[84][227], Harray[85][227], Harray[86][227], Harray[87][227], Harray[88][227], Harray[89][227], Harray[90][227], Harray[91][227], Harray[92][227], Harray[93][227], Harray[94][227], Harray[95][227], Harray[96][227], Harray[97][227], Harray[98][227], Harray[99][227], Harray[100][227], Harray[101][227], Harray[102][227], Harray[103][227], Harray[104][227], Harray[105][227], Harray[106][227], Harray[107][227], Harray[108][227], Harray[109][227], Harray[110][227], Harray[111][227], Harray[112][227], Harray[113][227], Harray[114][227], Harray[115][227], Harray[116][227], Harray[117][227], Harray[118][227], Harray[119][227], Harray[120][227], Harray[121][227], Harray[122][227], Harray[123][227], Harray[124][227], Harray[125][227], Harray[126][227], Harray[127][227]};
assign h_col_228 = {Harray[0][228], Harray[1][228], Harray[2][228], Harray[3][228], Harray[4][228], Harray[5][228], Harray[6][228], Harray[7][228], Harray[8][228], Harray[9][228], Harray[10][228], Harray[11][228], Harray[12][228], Harray[13][228], Harray[14][228], Harray[15][228], Harray[16][228], Harray[17][228], Harray[18][228], Harray[19][228], Harray[20][228], Harray[21][228], Harray[22][228], Harray[23][228], Harray[24][228], Harray[25][228], Harray[26][228], Harray[27][228], Harray[28][228], Harray[29][228], Harray[30][228], Harray[31][228], Harray[32][228], Harray[33][228], Harray[34][228], Harray[35][228], Harray[36][228], Harray[37][228], Harray[38][228], Harray[39][228], Harray[40][228], Harray[41][228], Harray[42][228], Harray[43][228], Harray[44][228], Harray[45][228], Harray[46][228], Harray[47][228], Harray[48][228], Harray[49][228], Harray[50][228], Harray[51][228], Harray[52][228], Harray[53][228], Harray[54][228], Harray[55][228], Harray[56][228], Harray[57][228], Harray[58][228], Harray[59][228], Harray[60][228], Harray[61][228], Harray[62][228], Harray[63][228], Harray[64][228], Harray[65][228], Harray[66][228], Harray[67][228], Harray[68][228], Harray[69][228], Harray[70][228], Harray[71][228], Harray[72][228], Harray[73][228], Harray[74][228], Harray[75][228], Harray[76][228], Harray[77][228], Harray[78][228], Harray[79][228], Harray[80][228], Harray[81][228], Harray[82][228], Harray[83][228], Harray[84][228], Harray[85][228], Harray[86][228], Harray[87][228], Harray[88][228], Harray[89][228], Harray[90][228], Harray[91][228], Harray[92][228], Harray[93][228], Harray[94][228], Harray[95][228], Harray[96][228], Harray[97][228], Harray[98][228], Harray[99][228], Harray[100][228], Harray[101][228], Harray[102][228], Harray[103][228], Harray[104][228], Harray[105][228], Harray[106][228], Harray[107][228], Harray[108][228], Harray[109][228], Harray[110][228], Harray[111][228], Harray[112][228], Harray[113][228], Harray[114][228], Harray[115][228], Harray[116][228], Harray[117][228], Harray[118][228], Harray[119][228], Harray[120][228], Harray[121][228], Harray[122][228], Harray[123][228], Harray[124][228], Harray[125][228], Harray[126][228], Harray[127][228]};
assign h_col_229 = {Harray[0][229], Harray[1][229], Harray[2][229], Harray[3][229], Harray[4][229], Harray[5][229], Harray[6][229], Harray[7][229], Harray[8][229], Harray[9][229], Harray[10][229], Harray[11][229], Harray[12][229], Harray[13][229], Harray[14][229], Harray[15][229], Harray[16][229], Harray[17][229], Harray[18][229], Harray[19][229], Harray[20][229], Harray[21][229], Harray[22][229], Harray[23][229], Harray[24][229], Harray[25][229], Harray[26][229], Harray[27][229], Harray[28][229], Harray[29][229], Harray[30][229], Harray[31][229], Harray[32][229], Harray[33][229], Harray[34][229], Harray[35][229], Harray[36][229], Harray[37][229], Harray[38][229], Harray[39][229], Harray[40][229], Harray[41][229], Harray[42][229], Harray[43][229], Harray[44][229], Harray[45][229], Harray[46][229], Harray[47][229], Harray[48][229], Harray[49][229], Harray[50][229], Harray[51][229], Harray[52][229], Harray[53][229], Harray[54][229], Harray[55][229], Harray[56][229], Harray[57][229], Harray[58][229], Harray[59][229], Harray[60][229], Harray[61][229], Harray[62][229], Harray[63][229], Harray[64][229], Harray[65][229], Harray[66][229], Harray[67][229], Harray[68][229], Harray[69][229], Harray[70][229], Harray[71][229], Harray[72][229], Harray[73][229], Harray[74][229], Harray[75][229], Harray[76][229], Harray[77][229], Harray[78][229], Harray[79][229], Harray[80][229], Harray[81][229], Harray[82][229], Harray[83][229], Harray[84][229], Harray[85][229], Harray[86][229], Harray[87][229], Harray[88][229], Harray[89][229], Harray[90][229], Harray[91][229], Harray[92][229], Harray[93][229], Harray[94][229], Harray[95][229], Harray[96][229], Harray[97][229], Harray[98][229], Harray[99][229], Harray[100][229], Harray[101][229], Harray[102][229], Harray[103][229], Harray[104][229], Harray[105][229], Harray[106][229], Harray[107][229], Harray[108][229], Harray[109][229], Harray[110][229], Harray[111][229], Harray[112][229], Harray[113][229], Harray[114][229], Harray[115][229], Harray[116][229], Harray[117][229], Harray[118][229], Harray[119][229], Harray[120][229], Harray[121][229], Harray[122][229], Harray[123][229], Harray[124][229], Harray[125][229], Harray[126][229], Harray[127][229]};
assign h_col_230 = {Harray[0][230], Harray[1][230], Harray[2][230], Harray[3][230], Harray[4][230], Harray[5][230], Harray[6][230], Harray[7][230], Harray[8][230], Harray[9][230], Harray[10][230], Harray[11][230], Harray[12][230], Harray[13][230], Harray[14][230], Harray[15][230], Harray[16][230], Harray[17][230], Harray[18][230], Harray[19][230], Harray[20][230], Harray[21][230], Harray[22][230], Harray[23][230], Harray[24][230], Harray[25][230], Harray[26][230], Harray[27][230], Harray[28][230], Harray[29][230], Harray[30][230], Harray[31][230], Harray[32][230], Harray[33][230], Harray[34][230], Harray[35][230], Harray[36][230], Harray[37][230], Harray[38][230], Harray[39][230], Harray[40][230], Harray[41][230], Harray[42][230], Harray[43][230], Harray[44][230], Harray[45][230], Harray[46][230], Harray[47][230], Harray[48][230], Harray[49][230], Harray[50][230], Harray[51][230], Harray[52][230], Harray[53][230], Harray[54][230], Harray[55][230], Harray[56][230], Harray[57][230], Harray[58][230], Harray[59][230], Harray[60][230], Harray[61][230], Harray[62][230], Harray[63][230], Harray[64][230], Harray[65][230], Harray[66][230], Harray[67][230], Harray[68][230], Harray[69][230], Harray[70][230], Harray[71][230], Harray[72][230], Harray[73][230], Harray[74][230], Harray[75][230], Harray[76][230], Harray[77][230], Harray[78][230], Harray[79][230], Harray[80][230], Harray[81][230], Harray[82][230], Harray[83][230], Harray[84][230], Harray[85][230], Harray[86][230], Harray[87][230], Harray[88][230], Harray[89][230], Harray[90][230], Harray[91][230], Harray[92][230], Harray[93][230], Harray[94][230], Harray[95][230], Harray[96][230], Harray[97][230], Harray[98][230], Harray[99][230], Harray[100][230], Harray[101][230], Harray[102][230], Harray[103][230], Harray[104][230], Harray[105][230], Harray[106][230], Harray[107][230], Harray[108][230], Harray[109][230], Harray[110][230], Harray[111][230], Harray[112][230], Harray[113][230], Harray[114][230], Harray[115][230], Harray[116][230], Harray[117][230], Harray[118][230], Harray[119][230], Harray[120][230], Harray[121][230], Harray[122][230], Harray[123][230], Harray[124][230], Harray[125][230], Harray[126][230], Harray[127][230]};
assign h_col_231 = {Harray[0][231], Harray[1][231], Harray[2][231], Harray[3][231], Harray[4][231], Harray[5][231], Harray[6][231], Harray[7][231], Harray[8][231], Harray[9][231], Harray[10][231], Harray[11][231], Harray[12][231], Harray[13][231], Harray[14][231], Harray[15][231], Harray[16][231], Harray[17][231], Harray[18][231], Harray[19][231], Harray[20][231], Harray[21][231], Harray[22][231], Harray[23][231], Harray[24][231], Harray[25][231], Harray[26][231], Harray[27][231], Harray[28][231], Harray[29][231], Harray[30][231], Harray[31][231], Harray[32][231], Harray[33][231], Harray[34][231], Harray[35][231], Harray[36][231], Harray[37][231], Harray[38][231], Harray[39][231], Harray[40][231], Harray[41][231], Harray[42][231], Harray[43][231], Harray[44][231], Harray[45][231], Harray[46][231], Harray[47][231], Harray[48][231], Harray[49][231], Harray[50][231], Harray[51][231], Harray[52][231], Harray[53][231], Harray[54][231], Harray[55][231], Harray[56][231], Harray[57][231], Harray[58][231], Harray[59][231], Harray[60][231], Harray[61][231], Harray[62][231], Harray[63][231], Harray[64][231], Harray[65][231], Harray[66][231], Harray[67][231], Harray[68][231], Harray[69][231], Harray[70][231], Harray[71][231], Harray[72][231], Harray[73][231], Harray[74][231], Harray[75][231], Harray[76][231], Harray[77][231], Harray[78][231], Harray[79][231], Harray[80][231], Harray[81][231], Harray[82][231], Harray[83][231], Harray[84][231], Harray[85][231], Harray[86][231], Harray[87][231], Harray[88][231], Harray[89][231], Harray[90][231], Harray[91][231], Harray[92][231], Harray[93][231], Harray[94][231], Harray[95][231], Harray[96][231], Harray[97][231], Harray[98][231], Harray[99][231], Harray[100][231], Harray[101][231], Harray[102][231], Harray[103][231], Harray[104][231], Harray[105][231], Harray[106][231], Harray[107][231], Harray[108][231], Harray[109][231], Harray[110][231], Harray[111][231], Harray[112][231], Harray[113][231], Harray[114][231], Harray[115][231], Harray[116][231], Harray[117][231], Harray[118][231], Harray[119][231], Harray[120][231], Harray[121][231], Harray[122][231], Harray[123][231], Harray[124][231], Harray[125][231], Harray[126][231], Harray[127][231]};
assign h_col_232 = {Harray[0][232], Harray[1][232], Harray[2][232], Harray[3][232], Harray[4][232], Harray[5][232], Harray[6][232], Harray[7][232], Harray[8][232], Harray[9][232], Harray[10][232], Harray[11][232], Harray[12][232], Harray[13][232], Harray[14][232], Harray[15][232], Harray[16][232], Harray[17][232], Harray[18][232], Harray[19][232], Harray[20][232], Harray[21][232], Harray[22][232], Harray[23][232], Harray[24][232], Harray[25][232], Harray[26][232], Harray[27][232], Harray[28][232], Harray[29][232], Harray[30][232], Harray[31][232], Harray[32][232], Harray[33][232], Harray[34][232], Harray[35][232], Harray[36][232], Harray[37][232], Harray[38][232], Harray[39][232], Harray[40][232], Harray[41][232], Harray[42][232], Harray[43][232], Harray[44][232], Harray[45][232], Harray[46][232], Harray[47][232], Harray[48][232], Harray[49][232], Harray[50][232], Harray[51][232], Harray[52][232], Harray[53][232], Harray[54][232], Harray[55][232], Harray[56][232], Harray[57][232], Harray[58][232], Harray[59][232], Harray[60][232], Harray[61][232], Harray[62][232], Harray[63][232], Harray[64][232], Harray[65][232], Harray[66][232], Harray[67][232], Harray[68][232], Harray[69][232], Harray[70][232], Harray[71][232], Harray[72][232], Harray[73][232], Harray[74][232], Harray[75][232], Harray[76][232], Harray[77][232], Harray[78][232], Harray[79][232], Harray[80][232], Harray[81][232], Harray[82][232], Harray[83][232], Harray[84][232], Harray[85][232], Harray[86][232], Harray[87][232], Harray[88][232], Harray[89][232], Harray[90][232], Harray[91][232], Harray[92][232], Harray[93][232], Harray[94][232], Harray[95][232], Harray[96][232], Harray[97][232], Harray[98][232], Harray[99][232], Harray[100][232], Harray[101][232], Harray[102][232], Harray[103][232], Harray[104][232], Harray[105][232], Harray[106][232], Harray[107][232], Harray[108][232], Harray[109][232], Harray[110][232], Harray[111][232], Harray[112][232], Harray[113][232], Harray[114][232], Harray[115][232], Harray[116][232], Harray[117][232], Harray[118][232], Harray[119][232], Harray[120][232], Harray[121][232], Harray[122][232], Harray[123][232], Harray[124][232], Harray[125][232], Harray[126][232], Harray[127][232]};
assign h_col_233 = {Harray[0][233], Harray[1][233], Harray[2][233], Harray[3][233], Harray[4][233], Harray[5][233], Harray[6][233], Harray[7][233], Harray[8][233], Harray[9][233], Harray[10][233], Harray[11][233], Harray[12][233], Harray[13][233], Harray[14][233], Harray[15][233], Harray[16][233], Harray[17][233], Harray[18][233], Harray[19][233], Harray[20][233], Harray[21][233], Harray[22][233], Harray[23][233], Harray[24][233], Harray[25][233], Harray[26][233], Harray[27][233], Harray[28][233], Harray[29][233], Harray[30][233], Harray[31][233], Harray[32][233], Harray[33][233], Harray[34][233], Harray[35][233], Harray[36][233], Harray[37][233], Harray[38][233], Harray[39][233], Harray[40][233], Harray[41][233], Harray[42][233], Harray[43][233], Harray[44][233], Harray[45][233], Harray[46][233], Harray[47][233], Harray[48][233], Harray[49][233], Harray[50][233], Harray[51][233], Harray[52][233], Harray[53][233], Harray[54][233], Harray[55][233], Harray[56][233], Harray[57][233], Harray[58][233], Harray[59][233], Harray[60][233], Harray[61][233], Harray[62][233], Harray[63][233], Harray[64][233], Harray[65][233], Harray[66][233], Harray[67][233], Harray[68][233], Harray[69][233], Harray[70][233], Harray[71][233], Harray[72][233], Harray[73][233], Harray[74][233], Harray[75][233], Harray[76][233], Harray[77][233], Harray[78][233], Harray[79][233], Harray[80][233], Harray[81][233], Harray[82][233], Harray[83][233], Harray[84][233], Harray[85][233], Harray[86][233], Harray[87][233], Harray[88][233], Harray[89][233], Harray[90][233], Harray[91][233], Harray[92][233], Harray[93][233], Harray[94][233], Harray[95][233], Harray[96][233], Harray[97][233], Harray[98][233], Harray[99][233], Harray[100][233], Harray[101][233], Harray[102][233], Harray[103][233], Harray[104][233], Harray[105][233], Harray[106][233], Harray[107][233], Harray[108][233], Harray[109][233], Harray[110][233], Harray[111][233], Harray[112][233], Harray[113][233], Harray[114][233], Harray[115][233], Harray[116][233], Harray[117][233], Harray[118][233], Harray[119][233], Harray[120][233], Harray[121][233], Harray[122][233], Harray[123][233], Harray[124][233], Harray[125][233], Harray[126][233], Harray[127][233]};
assign h_col_234 = {Harray[0][234], Harray[1][234], Harray[2][234], Harray[3][234], Harray[4][234], Harray[5][234], Harray[6][234], Harray[7][234], Harray[8][234], Harray[9][234], Harray[10][234], Harray[11][234], Harray[12][234], Harray[13][234], Harray[14][234], Harray[15][234], Harray[16][234], Harray[17][234], Harray[18][234], Harray[19][234], Harray[20][234], Harray[21][234], Harray[22][234], Harray[23][234], Harray[24][234], Harray[25][234], Harray[26][234], Harray[27][234], Harray[28][234], Harray[29][234], Harray[30][234], Harray[31][234], Harray[32][234], Harray[33][234], Harray[34][234], Harray[35][234], Harray[36][234], Harray[37][234], Harray[38][234], Harray[39][234], Harray[40][234], Harray[41][234], Harray[42][234], Harray[43][234], Harray[44][234], Harray[45][234], Harray[46][234], Harray[47][234], Harray[48][234], Harray[49][234], Harray[50][234], Harray[51][234], Harray[52][234], Harray[53][234], Harray[54][234], Harray[55][234], Harray[56][234], Harray[57][234], Harray[58][234], Harray[59][234], Harray[60][234], Harray[61][234], Harray[62][234], Harray[63][234], Harray[64][234], Harray[65][234], Harray[66][234], Harray[67][234], Harray[68][234], Harray[69][234], Harray[70][234], Harray[71][234], Harray[72][234], Harray[73][234], Harray[74][234], Harray[75][234], Harray[76][234], Harray[77][234], Harray[78][234], Harray[79][234], Harray[80][234], Harray[81][234], Harray[82][234], Harray[83][234], Harray[84][234], Harray[85][234], Harray[86][234], Harray[87][234], Harray[88][234], Harray[89][234], Harray[90][234], Harray[91][234], Harray[92][234], Harray[93][234], Harray[94][234], Harray[95][234], Harray[96][234], Harray[97][234], Harray[98][234], Harray[99][234], Harray[100][234], Harray[101][234], Harray[102][234], Harray[103][234], Harray[104][234], Harray[105][234], Harray[106][234], Harray[107][234], Harray[108][234], Harray[109][234], Harray[110][234], Harray[111][234], Harray[112][234], Harray[113][234], Harray[114][234], Harray[115][234], Harray[116][234], Harray[117][234], Harray[118][234], Harray[119][234], Harray[120][234], Harray[121][234], Harray[122][234], Harray[123][234], Harray[124][234], Harray[125][234], Harray[126][234], Harray[127][234]};
assign h_col_235 = {Harray[0][235], Harray[1][235], Harray[2][235], Harray[3][235], Harray[4][235], Harray[5][235], Harray[6][235], Harray[7][235], Harray[8][235], Harray[9][235], Harray[10][235], Harray[11][235], Harray[12][235], Harray[13][235], Harray[14][235], Harray[15][235], Harray[16][235], Harray[17][235], Harray[18][235], Harray[19][235], Harray[20][235], Harray[21][235], Harray[22][235], Harray[23][235], Harray[24][235], Harray[25][235], Harray[26][235], Harray[27][235], Harray[28][235], Harray[29][235], Harray[30][235], Harray[31][235], Harray[32][235], Harray[33][235], Harray[34][235], Harray[35][235], Harray[36][235], Harray[37][235], Harray[38][235], Harray[39][235], Harray[40][235], Harray[41][235], Harray[42][235], Harray[43][235], Harray[44][235], Harray[45][235], Harray[46][235], Harray[47][235], Harray[48][235], Harray[49][235], Harray[50][235], Harray[51][235], Harray[52][235], Harray[53][235], Harray[54][235], Harray[55][235], Harray[56][235], Harray[57][235], Harray[58][235], Harray[59][235], Harray[60][235], Harray[61][235], Harray[62][235], Harray[63][235], Harray[64][235], Harray[65][235], Harray[66][235], Harray[67][235], Harray[68][235], Harray[69][235], Harray[70][235], Harray[71][235], Harray[72][235], Harray[73][235], Harray[74][235], Harray[75][235], Harray[76][235], Harray[77][235], Harray[78][235], Harray[79][235], Harray[80][235], Harray[81][235], Harray[82][235], Harray[83][235], Harray[84][235], Harray[85][235], Harray[86][235], Harray[87][235], Harray[88][235], Harray[89][235], Harray[90][235], Harray[91][235], Harray[92][235], Harray[93][235], Harray[94][235], Harray[95][235], Harray[96][235], Harray[97][235], Harray[98][235], Harray[99][235], Harray[100][235], Harray[101][235], Harray[102][235], Harray[103][235], Harray[104][235], Harray[105][235], Harray[106][235], Harray[107][235], Harray[108][235], Harray[109][235], Harray[110][235], Harray[111][235], Harray[112][235], Harray[113][235], Harray[114][235], Harray[115][235], Harray[116][235], Harray[117][235], Harray[118][235], Harray[119][235], Harray[120][235], Harray[121][235], Harray[122][235], Harray[123][235], Harray[124][235], Harray[125][235], Harray[126][235], Harray[127][235]};
assign h_col_236 = {Harray[0][236], Harray[1][236], Harray[2][236], Harray[3][236], Harray[4][236], Harray[5][236], Harray[6][236], Harray[7][236], Harray[8][236], Harray[9][236], Harray[10][236], Harray[11][236], Harray[12][236], Harray[13][236], Harray[14][236], Harray[15][236], Harray[16][236], Harray[17][236], Harray[18][236], Harray[19][236], Harray[20][236], Harray[21][236], Harray[22][236], Harray[23][236], Harray[24][236], Harray[25][236], Harray[26][236], Harray[27][236], Harray[28][236], Harray[29][236], Harray[30][236], Harray[31][236], Harray[32][236], Harray[33][236], Harray[34][236], Harray[35][236], Harray[36][236], Harray[37][236], Harray[38][236], Harray[39][236], Harray[40][236], Harray[41][236], Harray[42][236], Harray[43][236], Harray[44][236], Harray[45][236], Harray[46][236], Harray[47][236], Harray[48][236], Harray[49][236], Harray[50][236], Harray[51][236], Harray[52][236], Harray[53][236], Harray[54][236], Harray[55][236], Harray[56][236], Harray[57][236], Harray[58][236], Harray[59][236], Harray[60][236], Harray[61][236], Harray[62][236], Harray[63][236], Harray[64][236], Harray[65][236], Harray[66][236], Harray[67][236], Harray[68][236], Harray[69][236], Harray[70][236], Harray[71][236], Harray[72][236], Harray[73][236], Harray[74][236], Harray[75][236], Harray[76][236], Harray[77][236], Harray[78][236], Harray[79][236], Harray[80][236], Harray[81][236], Harray[82][236], Harray[83][236], Harray[84][236], Harray[85][236], Harray[86][236], Harray[87][236], Harray[88][236], Harray[89][236], Harray[90][236], Harray[91][236], Harray[92][236], Harray[93][236], Harray[94][236], Harray[95][236], Harray[96][236], Harray[97][236], Harray[98][236], Harray[99][236], Harray[100][236], Harray[101][236], Harray[102][236], Harray[103][236], Harray[104][236], Harray[105][236], Harray[106][236], Harray[107][236], Harray[108][236], Harray[109][236], Harray[110][236], Harray[111][236], Harray[112][236], Harray[113][236], Harray[114][236], Harray[115][236], Harray[116][236], Harray[117][236], Harray[118][236], Harray[119][236], Harray[120][236], Harray[121][236], Harray[122][236], Harray[123][236], Harray[124][236], Harray[125][236], Harray[126][236], Harray[127][236]};
assign h_col_237 = {Harray[0][237], Harray[1][237], Harray[2][237], Harray[3][237], Harray[4][237], Harray[5][237], Harray[6][237], Harray[7][237], Harray[8][237], Harray[9][237], Harray[10][237], Harray[11][237], Harray[12][237], Harray[13][237], Harray[14][237], Harray[15][237], Harray[16][237], Harray[17][237], Harray[18][237], Harray[19][237], Harray[20][237], Harray[21][237], Harray[22][237], Harray[23][237], Harray[24][237], Harray[25][237], Harray[26][237], Harray[27][237], Harray[28][237], Harray[29][237], Harray[30][237], Harray[31][237], Harray[32][237], Harray[33][237], Harray[34][237], Harray[35][237], Harray[36][237], Harray[37][237], Harray[38][237], Harray[39][237], Harray[40][237], Harray[41][237], Harray[42][237], Harray[43][237], Harray[44][237], Harray[45][237], Harray[46][237], Harray[47][237], Harray[48][237], Harray[49][237], Harray[50][237], Harray[51][237], Harray[52][237], Harray[53][237], Harray[54][237], Harray[55][237], Harray[56][237], Harray[57][237], Harray[58][237], Harray[59][237], Harray[60][237], Harray[61][237], Harray[62][237], Harray[63][237], Harray[64][237], Harray[65][237], Harray[66][237], Harray[67][237], Harray[68][237], Harray[69][237], Harray[70][237], Harray[71][237], Harray[72][237], Harray[73][237], Harray[74][237], Harray[75][237], Harray[76][237], Harray[77][237], Harray[78][237], Harray[79][237], Harray[80][237], Harray[81][237], Harray[82][237], Harray[83][237], Harray[84][237], Harray[85][237], Harray[86][237], Harray[87][237], Harray[88][237], Harray[89][237], Harray[90][237], Harray[91][237], Harray[92][237], Harray[93][237], Harray[94][237], Harray[95][237], Harray[96][237], Harray[97][237], Harray[98][237], Harray[99][237], Harray[100][237], Harray[101][237], Harray[102][237], Harray[103][237], Harray[104][237], Harray[105][237], Harray[106][237], Harray[107][237], Harray[108][237], Harray[109][237], Harray[110][237], Harray[111][237], Harray[112][237], Harray[113][237], Harray[114][237], Harray[115][237], Harray[116][237], Harray[117][237], Harray[118][237], Harray[119][237], Harray[120][237], Harray[121][237], Harray[122][237], Harray[123][237], Harray[124][237], Harray[125][237], Harray[126][237], Harray[127][237]};
assign h_col_238 = {Harray[0][238], Harray[1][238], Harray[2][238], Harray[3][238], Harray[4][238], Harray[5][238], Harray[6][238], Harray[7][238], Harray[8][238], Harray[9][238], Harray[10][238], Harray[11][238], Harray[12][238], Harray[13][238], Harray[14][238], Harray[15][238], Harray[16][238], Harray[17][238], Harray[18][238], Harray[19][238], Harray[20][238], Harray[21][238], Harray[22][238], Harray[23][238], Harray[24][238], Harray[25][238], Harray[26][238], Harray[27][238], Harray[28][238], Harray[29][238], Harray[30][238], Harray[31][238], Harray[32][238], Harray[33][238], Harray[34][238], Harray[35][238], Harray[36][238], Harray[37][238], Harray[38][238], Harray[39][238], Harray[40][238], Harray[41][238], Harray[42][238], Harray[43][238], Harray[44][238], Harray[45][238], Harray[46][238], Harray[47][238], Harray[48][238], Harray[49][238], Harray[50][238], Harray[51][238], Harray[52][238], Harray[53][238], Harray[54][238], Harray[55][238], Harray[56][238], Harray[57][238], Harray[58][238], Harray[59][238], Harray[60][238], Harray[61][238], Harray[62][238], Harray[63][238], Harray[64][238], Harray[65][238], Harray[66][238], Harray[67][238], Harray[68][238], Harray[69][238], Harray[70][238], Harray[71][238], Harray[72][238], Harray[73][238], Harray[74][238], Harray[75][238], Harray[76][238], Harray[77][238], Harray[78][238], Harray[79][238], Harray[80][238], Harray[81][238], Harray[82][238], Harray[83][238], Harray[84][238], Harray[85][238], Harray[86][238], Harray[87][238], Harray[88][238], Harray[89][238], Harray[90][238], Harray[91][238], Harray[92][238], Harray[93][238], Harray[94][238], Harray[95][238], Harray[96][238], Harray[97][238], Harray[98][238], Harray[99][238], Harray[100][238], Harray[101][238], Harray[102][238], Harray[103][238], Harray[104][238], Harray[105][238], Harray[106][238], Harray[107][238], Harray[108][238], Harray[109][238], Harray[110][238], Harray[111][238], Harray[112][238], Harray[113][238], Harray[114][238], Harray[115][238], Harray[116][238], Harray[117][238], Harray[118][238], Harray[119][238], Harray[120][238], Harray[121][238], Harray[122][238], Harray[123][238], Harray[124][238], Harray[125][238], Harray[126][238], Harray[127][238]};
assign h_col_239 = {Harray[0][239], Harray[1][239], Harray[2][239], Harray[3][239], Harray[4][239], Harray[5][239], Harray[6][239], Harray[7][239], Harray[8][239], Harray[9][239], Harray[10][239], Harray[11][239], Harray[12][239], Harray[13][239], Harray[14][239], Harray[15][239], Harray[16][239], Harray[17][239], Harray[18][239], Harray[19][239], Harray[20][239], Harray[21][239], Harray[22][239], Harray[23][239], Harray[24][239], Harray[25][239], Harray[26][239], Harray[27][239], Harray[28][239], Harray[29][239], Harray[30][239], Harray[31][239], Harray[32][239], Harray[33][239], Harray[34][239], Harray[35][239], Harray[36][239], Harray[37][239], Harray[38][239], Harray[39][239], Harray[40][239], Harray[41][239], Harray[42][239], Harray[43][239], Harray[44][239], Harray[45][239], Harray[46][239], Harray[47][239], Harray[48][239], Harray[49][239], Harray[50][239], Harray[51][239], Harray[52][239], Harray[53][239], Harray[54][239], Harray[55][239], Harray[56][239], Harray[57][239], Harray[58][239], Harray[59][239], Harray[60][239], Harray[61][239], Harray[62][239], Harray[63][239], Harray[64][239], Harray[65][239], Harray[66][239], Harray[67][239], Harray[68][239], Harray[69][239], Harray[70][239], Harray[71][239], Harray[72][239], Harray[73][239], Harray[74][239], Harray[75][239], Harray[76][239], Harray[77][239], Harray[78][239], Harray[79][239], Harray[80][239], Harray[81][239], Harray[82][239], Harray[83][239], Harray[84][239], Harray[85][239], Harray[86][239], Harray[87][239], Harray[88][239], Harray[89][239], Harray[90][239], Harray[91][239], Harray[92][239], Harray[93][239], Harray[94][239], Harray[95][239], Harray[96][239], Harray[97][239], Harray[98][239], Harray[99][239], Harray[100][239], Harray[101][239], Harray[102][239], Harray[103][239], Harray[104][239], Harray[105][239], Harray[106][239], Harray[107][239], Harray[108][239], Harray[109][239], Harray[110][239], Harray[111][239], Harray[112][239], Harray[113][239], Harray[114][239], Harray[115][239], Harray[116][239], Harray[117][239], Harray[118][239], Harray[119][239], Harray[120][239], Harray[121][239], Harray[122][239], Harray[123][239], Harray[124][239], Harray[125][239], Harray[126][239], Harray[127][239]};
assign h_col_240 = {Harray[0][240], Harray[1][240], Harray[2][240], Harray[3][240], Harray[4][240], Harray[5][240], Harray[6][240], Harray[7][240], Harray[8][240], Harray[9][240], Harray[10][240], Harray[11][240], Harray[12][240], Harray[13][240], Harray[14][240], Harray[15][240], Harray[16][240], Harray[17][240], Harray[18][240], Harray[19][240], Harray[20][240], Harray[21][240], Harray[22][240], Harray[23][240], Harray[24][240], Harray[25][240], Harray[26][240], Harray[27][240], Harray[28][240], Harray[29][240], Harray[30][240], Harray[31][240], Harray[32][240], Harray[33][240], Harray[34][240], Harray[35][240], Harray[36][240], Harray[37][240], Harray[38][240], Harray[39][240], Harray[40][240], Harray[41][240], Harray[42][240], Harray[43][240], Harray[44][240], Harray[45][240], Harray[46][240], Harray[47][240], Harray[48][240], Harray[49][240], Harray[50][240], Harray[51][240], Harray[52][240], Harray[53][240], Harray[54][240], Harray[55][240], Harray[56][240], Harray[57][240], Harray[58][240], Harray[59][240], Harray[60][240], Harray[61][240], Harray[62][240], Harray[63][240], Harray[64][240], Harray[65][240], Harray[66][240], Harray[67][240], Harray[68][240], Harray[69][240], Harray[70][240], Harray[71][240], Harray[72][240], Harray[73][240], Harray[74][240], Harray[75][240], Harray[76][240], Harray[77][240], Harray[78][240], Harray[79][240], Harray[80][240], Harray[81][240], Harray[82][240], Harray[83][240], Harray[84][240], Harray[85][240], Harray[86][240], Harray[87][240], Harray[88][240], Harray[89][240], Harray[90][240], Harray[91][240], Harray[92][240], Harray[93][240], Harray[94][240], Harray[95][240], Harray[96][240], Harray[97][240], Harray[98][240], Harray[99][240], Harray[100][240], Harray[101][240], Harray[102][240], Harray[103][240], Harray[104][240], Harray[105][240], Harray[106][240], Harray[107][240], Harray[108][240], Harray[109][240], Harray[110][240], Harray[111][240], Harray[112][240], Harray[113][240], Harray[114][240], Harray[115][240], Harray[116][240], Harray[117][240], Harray[118][240], Harray[119][240], Harray[120][240], Harray[121][240], Harray[122][240], Harray[123][240], Harray[124][240], Harray[125][240], Harray[126][240], Harray[127][240]};
assign h_col_241 = {Harray[0][241], Harray[1][241], Harray[2][241], Harray[3][241], Harray[4][241], Harray[5][241], Harray[6][241], Harray[7][241], Harray[8][241], Harray[9][241], Harray[10][241], Harray[11][241], Harray[12][241], Harray[13][241], Harray[14][241], Harray[15][241], Harray[16][241], Harray[17][241], Harray[18][241], Harray[19][241], Harray[20][241], Harray[21][241], Harray[22][241], Harray[23][241], Harray[24][241], Harray[25][241], Harray[26][241], Harray[27][241], Harray[28][241], Harray[29][241], Harray[30][241], Harray[31][241], Harray[32][241], Harray[33][241], Harray[34][241], Harray[35][241], Harray[36][241], Harray[37][241], Harray[38][241], Harray[39][241], Harray[40][241], Harray[41][241], Harray[42][241], Harray[43][241], Harray[44][241], Harray[45][241], Harray[46][241], Harray[47][241], Harray[48][241], Harray[49][241], Harray[50][241], Harray[51][241], Harray[52][241], Harray[53][241], Harray[54][241], Harray[55][241], Harray[56][241], Harray[57][241], Harray[58][241], Harray[59][241], Harray[60][241], Harray[61][241], Harray[62][241], Harray[63][241], Harray[64][241], Harray[65][241], Harray[66][241], Harray[67][241], Harray[68][241], Harray[69][241], Harray[70][241], Harray[71][241], Harray[72][241], Harray[73][241], Harray[74][241], Harray[75][241], Harray[76][241], Harray[77][241], Harray[78][241], Harray[79][241], Harray[80][241], Harray[81][241], Harray[82][241], Harray[83][241], Harray[84][241], Harray[85][241], Harray[86][241], Harray[87][241], Harray[88][241], Harray[89][241], Harray[90][241], Harray[91][241], Harray[92][241], Harray[93][241], Harray[94][241], Harray[95][241], Harray[96][241], Harray[97][241], Harray[98][241], Harray[99][241], Harray[100][241], Harray[101][241], Harray[102][241], Harray[103][241], Harray[104][241], Harray[105][241], Harray[106][241], Harray[107][241], Harray[108][241], Harray[109][241], Harray[110][241], Harray[111][241], Harray[112][241], Harray[113][241], Harray[114][241], Harray[115][241], Harray[116][241], Harray[117][241], Harray[118][241], Harray[119][241], Harray[120][241], Harray[121][241], Harray[122][241], Harray[123][241], Harray[124][241], Harray[125][241], Harray[126][241], Harray[127][241]};
assign h_col_242 = {Harray[0][242], Harray[1][242], Harray[2][242], Harray[3][242], Harray[4][242], Harray[5][242], Harray[6][242], Harray[7][242], Harray[8][242], Harray[9][242], Harray[10][242], Harray[11][242], Harray[12][242], Harray[13][242], Harray[14][242], Harray[15][242], Harray[16][242], Harray[17][242], Harray[18][242], Harray[19][242], Harray[20][242], Harray[21][242], Harray[22][242], Harray[23][242], Harray[24][242], Harray[25][242], Harray[26][242], Harray[27][242], Harray[28][242], Harray[29][242], Harray[30][242], Harray[31][242], Harray[32][242], Harray[33][242], Harray[34][242], Harray[35][242], Harray[36][242], Harray[37][242], Harray[38][242], Harray[39][242], Harray[40][242], Harray[41][242], Harray[42][242], Harray[43][242], Harray[44][242], Harray[45][242], Harray[46][242], Harray[47][242], Harray[48][242], Harray[49][242], Harray[50][242], Harray[51][242], Harray[52][242], Harray[53][242], Harray[54][242], Harray[55][242], Harray[56][242], Harray[57][242], Harray[58][242], Harray[59][242], Harray[60][242], Harray[61][242], Harray[62][242], Harray[63][242], Harray[64][242], Harray[65][242], Harray[66][242], Harray[67][242], Harray[68][242], Harray[69][242], Harray[70][242], Harray[71][242], Harray[72][242], Harray[73][242], Harray[74][242], Harray[75][242], Harray[76][242], Harray[77][242], Harray[78][242], Harray[79][242], Harray[80][242], Harray[81][242], Harray[82][242], Harray[83][242], Harray[84][242], Harray[85][242], Harray[86][242], Harray[87][242], Harray[88][242], Harray[89][242], Harray[90][242], Harray[91][242], Harray[92][242], Harray[93][242], Harray[94][242], Harray[95][242], Harray[96][242], Harray[97][242], Harray[98][242], Harray[99][242], Harray[100][242], Harray[101][242], Harray[102][242], Harray[103][242], Harray[104][242], Harray[105][242], Harray[106][242], Harray[107][242], Harray[108][242], Harray[109][242], Harray[110][242], Harray[111][242], Harray[112][242], Harray[113][242], Harray[114][242], Harray[115][242], Harray[116][242], Harray[117][242], Harray[118][242], Harray[119][242], Harray[120][242], Harray[121][242], Harray[122][242], Harray[123][242], Harray[124][242], Harray[125][242], Harray[126][242], Harray[127][242]};
assign h_col_243 = {Harray[0][243], Harray[1][243], Harray[2][243], Harray[3][243], Harray[4][243], Harray[5][243], Harray[6][243], Harray[7][243], Harray[8][243], Harray[9][243], Harray[10][243], Harray[11][243], Harray[12][243], Harray[13][243], Harray[14][243], Harray[15][243], Harray[16][243], Harray[17][243], Harray[18][243], Harray[19][243], Harray[20][243], Harray[21][243], Harray[22][243], Harray[23][243], Harray[24][243], Harray[25][243], Harray[26][243], Harray[27][243], Harray[28][243], Harray[29][243], Harray[30][243], Harray[31][243], Harray[32][243], Harray[33][243], Harray[34][243], Harray[35][243], Harray[36][243], Harray[37][243], Harray[38][243], Harray[39][243], Harray[40][243], Harray[41][243], Harray[42][243], Harray[43][243], Harray[44][243], Harray[45][243], Harray[46][243], Harray[47][243], Harray[48][243], Harray[49][243], Harray[50][243], Harray[51][243], Harray[52][243], Harray[53][243], Harray[54][243], Harray[55][243], Harray[56][243], Harray[57][243], Harray[58][243], Harray[59][243], Harray[60][243], Harray[61][243], Harray[62][243], Harray[63][243], Harray[64][243], Harray[65][243], Harray[66][243], Harray[67][243], Harray[68][243], Harray[69][243], Harray[70][243], Harray[71][243], Harray[72][243], Harray[73][243], Harray[74][243], Harray[75][243], Harray[76][243], Harray[77][243], Harray[78][243], Harray[79][243], Harray[80][243], Harray[81][243], Harray[82][243], Harray[83][243], Harray[84][243], Harray[85][243], Harray[86][243], Harray[87][243], Harray[88][243], Harray[89][243], Harray[90][243], Harray[91][243], Harray[92][243], Harray[93][243], Harray[94][243], Harray[95][243], Harray[96][243], Harray[97][243], Harray[98][243], Harray[99][243], Harray[100][243], Harray[101][243], Harray[102][243], Harray[103][243], Harray[104][243], Harray[105][243], Harray[106][243], Harray[107][243], Harray[108][243], Harray[109][243], Harray[110][243], Harray[111][243], Harray[112][243], Harray[113][243], Harray[114][243], Harray[115][243], Harray[116][243], Harray[117][243], Harray[118][243], Harray[119][243], Harray[120][243], Harray[121][243], Harray[122][243], Harray[123][243], Harray[124][243], Harray[125][243], Harray[126][243], Harray[127][243]};
assign h_col_244 = {Harray[0][244], Harray[1][244], Harray[2][244], Harray[3][244], Harray[4][244], Harray[5][244], Harray[6][244], Harray[7][244], Harray[8][244], Harray[9][244], Harray[10][244], Harray[11][244], Harray[12][244], Harray[13][244], Harray[14][244], Harray[15][244], Harray[16][244], Harray[17][244], Harray[18][244], Harray[19][244], Harray[20][244], Harray[21][244], Harray[22][244], Harray[23][244], Harray[24][244], Harray[25][244], Harray[26][244], Harray[27][244], Harray[28][244], Harray[29][244], Harray[30][244], Harray[31][244], Harray[32][244], Harray[33][244], Harray[34][244], Harray[35][244], Harray[36][244], Harray[37][244], Harray[38][244], Harray[39][244], Harray[40][244], Harray[41][244], Harray[42][244], Harray[43][244], Harray[44][244], Harray[45][244], Harray[46][244], Harray[47][244], Harray[48][244], Harray[49][244], Harray[50][244], Harray[51][244], Harray[52][244], Harray[53][244], Harray[54][244], Harray[55][244], Harray[56][244], Harray[57][244], Harray[58][244], Harray[59][244], Harray[60][244], Harray[61][244], Harray[62][244], Harray[63][244], Harray[64][244], Harray[65][244], Harray[66][244], Harray[67][244], Harray[68][244], Harray[69][244], Harray[70][244], Harray[71][244], Harray[72][244], Harray[73][244], Harray[74][244], Harray[75][244], Harray[76][244], Harray[77][244], Harray[78][244], Harray[79][244], Harray[80][244], Harray[81][244], Harray[82][244], Harray[83][244], Harray[84][244], Harray[85][244], Harray[86][244], Harray[87][244], Harray[88][244], Harray[89][244], Harray[90][244], Harray[91][244], Harray[92][244], Harray[93][244], Harray[94][244], Harray[95][244], Harray[96][244], Harray[97][244], Harray[98][244], Harray[99][244], Harray[100][244], Harray[101][244], Harray[102][244], Harray[103][244], Harray[104][244], Harray[105][244], Harray[106][244], Harray[107][244], Harray[108][244], Harray[109][244], Harray[110][244], Harray[111][244], Harray[112][244], Harray[113][244], Harray[114][244], Harray[115][244], Harray[116][244], Harray[117][244], Harray[118][244], Harray[119][244], Harray[120][244], Harray[121][244], Harray[122][244], Harray[123][244], Harray[124][244], Harray[125][244], Harray[126][244], Harray[127][244]};
assign h_col_245 = {Harray[0][245], Harray[1][245], Harray[2][245], Harray[3][245], Harray[4][245], Harray[5][245], Harray[6][245], Harray[7][245], Harray[8][245], Harray[9][245], Harray[10][245], Harray[11][245], Harray[12][245], Harray[13][245], Harray[14][245], Harray[15][245], Harray[16][245], Harray[17][245], Harray[18][245], Harray[19][245], Harray[20][245], Harray[21][245], Harray[22][245], Harray[23][245], Harray[24][245], Harray[25][245], Harray[26][245], Harray[27][245], Harray[28][245], Harray[29][245], Harray[30][245], Harray[31][245], Harray[32][245], Harray[33][245], Harray[34][245], Harray[35][245], Harray[36][245], Harray[37][245], Harray[38][245], Harray[39][245], Harray[40][245], Harray[41][245], Harray[42][245], Harray[43][245], Harray[44][245], Harray[45][245], Harray[46][245], Harray[47][245], Harray[48][245], Harray[49][245], Harray[50][245], Harray[51][245], Harray[52][245], Harray[53][245], Harray[54][245], Harray[55][245], Harray[56][245], Harray[57][245], Harray[58][245], Harray[59][245], Harray[60][245], Harray[61][245], Harray[62][245], Harray[63][245], Harray[64][245], Harray[65][245], Harray[66][245], Harray[67][245], Harray[68][245], Harray[69][245], Harray[70][245], Harray[71][245], Harray[72][245], Harray[73][245], Harray[74][245], Harray[75][245], Harray[76][245], Harray[77][245], Harray[78][245], Harray[79][245], Harray[80][245], Harray[81][245], Harray[82][245], Harray[83][245], Harray[84][245], Harray[85][245], Harray[86][245], Harray[87][245], Harray[88][245], Harray[89][245], Harray[90][245], Harray[91][245], Harray[92][245], Harray[93][245], Harray[94][245], Harray[95][245], Harray[96][245], Harray[97][245], Harray[98][245], Harray[99][245], Harray[100][245], Harray[101][245], Harray[102][245], Harray[103][245], Harray[104][245], Harray[105][245], Harray[106][245], Harray[107][245], Harray[108][245], Harray[109][245], Harray[110][245], Harray[111][245], Harray[112][245], Harray[113][245], Harray[114][245], Harray[115][245], Harray[116][245], Harray[117][245], Harray[118][245], Harray[119][245], Harray[120][245], Harray[121][245], Harray[122][245], Harray[123][245], Harray[124][245], Harray[125][245], Harray[126][245], Harray[127][245]};
assign h_col_246 = {Harray[0][246], Harray[1][246], Harray[2][246], Harray[3][246], Harray[4][246], Harray[5][246], Harray[6][246], Harray[7][246], Harray[8][246], Harray[9][246], Harray[10][246], Harray[11][246], Harray[12][246], Harray[13][246], Harray[14][246], Harray[15][246], Harray[16][246], Harray[17][246], Harray[18][246], Harray[19][246], Harray[20][246], Harray[21][246], Harray[22][246], Harray[23][246], Harray[24][246], Harray[25][246], Harray[26][246], Harray[27][246], Harray[28][246], Harray[29][246], Harray[30][246], Harray[31][246], Harray[32][246], Harray[33][246], Harray[34][246], Harray[35][246], Harray[36][246], Harray[37][246], Harray[38][246], Harray[39][246], Harray[40][246], Harray[41][246], Harray[42][246], Harray[43][246], Harray[44][246], Harray[45][246], Harray[46][246], Harray[47][246], Harray[48][246], Harray[49][246], Harray[50][246], Harray[51][246], Harray[52][246], Harray[53][246], Harray[54][246], Harray[55][246], Harray[56][246], Harray[57][246], Harray[58][246], Harray[59][246], Harray[60][246], Harray[61][246], Harray[62][246], Harray[63][246], Harray[64][246], Harray[65][246], Harray[66][246], Harray[67][246], Harray[68][246], Harray[69][246], Harray[70][246], Harray[71][246], Harray[72][246], Harray[73][246], Harray[74][246], Harray[75][246], Harray[76][246], Harray[77][246], Harray[78][246], Harray[79][246], Harray[80][246], Harray[81][246], Harray[82][246], Harray[83][246], Harray[84][246], Harray[85][246], Harray[86][246], Harray[87][246], Harray[88][246], Harray[89][246], Harray[90][246], Harray[91][246], Harray[92][246], Harray[93][246], Harray[94][246], Harray[95][246], Harray[96][246], Harray[97][246], Harray[98][246], Harray[99][246], Harray[100][246], Harray[101][246], Harray[102][246], Harray[103][246], Harray[104][246], Harray[105][246], Harray[106][246], Harray[107][246], Harray[108][246], Harray[109][246], Harray[110][246], Harray[111][246], Harray[112][246], Harray[113][246], Harray[114][246], Harray[115][246], Harray[116][246], Harray[117][246], Harray[118][246], Harray[119][246], Harray[120][246], Harray[121][246], Harray[122][246], Harray[123][246], Harray[124][246], Harray[125][246], Harray[126][246], Harray[127][246]};
assign h_col_247 = {Harray[0][247], Harray[1][247], Harray[2][247], Harray[3][247], Harray[4][247], Harray[5][247], Harray[6][247], Harray[7][247], Harray[8][247], Harray[9][247], Harray[10][247], Harray[11][247], Harray[12][247], Harray[13][247], Harray[14][247], Harray[15][247], Harray[16][247], Harray[17][247], Harray[18][247], Harray[19][247], Harray[20][247], Harray[21][247], Harray[22][247], Harray[23][247], Harray[24][247], Harray[25][247], Harray[26][247], Harray[27][247], Harray[28][247], Harray[29][247], Harray[30][247], Harray[31][247], Harray[32][247], Harray[33][247], Harray[34][247], Harray[35][247], Harray[36][247], Harray[37][247], Harray[38][247], Harray[39][247], Harray[40][247], Harray[41][247], Harray[42][247], Harray[43][247], Harray[44][247], Harray[45][247], Harray[46][247], Harray[47][247], Harray[48][247], Harray[49][247], Harray[50][247], Harray[51][247], Harray[52][247], Harray[53][247], Harray[54][247], Harray[55][247], Harray[56][247], Harray[57][247], Harray[58][247], Harray[59][247], Harray[60][247], Harray[61][247], Harray[62][247], Harray[63][247], Harray[64][247], Harray[65][247], Harray[66][247], Harray[67][247], Harray[68][247], Harray[69][247], Harray[70][247], Harray[71][247], Harray[72][247], Harray[73][247], Harray[74][247], Harray[75][247], Harray[76][247], Harray[77][247], Harray[78][247], Harray[79][247], Harray[80][247], Harray[81][247], Harray[82][247], Harray[83][247], Harray[84][247], Harray[85][247], Harray[86][247], Harray[87][247], Harray[88][247], Harray[89][247], Harray[90][247], Harray[91][247], Harray[92][247], Harray[93][247], Harray[94][247], Harray[95][247], Harray[96][247], Harray[97][247], Harray[98][247], Harray[99][247], Harray[100][247], Harray[101][247], Harray[102][247], Harray[103][247], Harray[104][247], Harray[105][247], Harray[106][247], Harray[107][247], Harray[108][247], Harray[109][247], Harray[110][247], Harray[111][247], Harray[112][247], Harray[113][247], Harray[114][247], Harray[115][247], Harray[116][247], Harray[117][247], Harray[118][247], Harray[119][247], Harray[120][247], Harray[121][247], Harray[122][247], Harray[123][247], Harray[124][247], Harray[125][247], Harray[126][247], Harray[127][247]};
assign h_col_248 = {Harray[0][248], Harray[1][248], Harray[2][248], Harray[3][248], Harray[4][248], Harray[5][248], Harray[6][248], Harray[7][248], Harray[8][248], Harray[9][248], Harray[10][248], Harray[11][248], Harray[12][248], Harray[13][248], Harray[14][248], Harray[15][248], Harray[16][248], Harray[17][248], Harray[18][248], Harray[19][248], Harray[20][248], Harray[21][248], Harray[22][248], Harray[23][248], Harray[24][248], Harray[25][248], Harray[26][248], Harray[27][248], Harray[28][248], Harray[29][248], Harray[30][248], Harray[31][248], Harray[32][248], Harray[33][248], Harray[34][248], Harray[35][248], Harray[36][248], Harray[37][248], Harray[38][248], Harray[39][248], Harray[40][248], Harray[41][248], Harray[42][248], Harray[43][248], Harray[44][248], Harray[45][248], Harray[46][248], Harray[47][248], Harray[48][248], Harray[49][248], Harray[50][248], Harray[51][248], Harray[52][248], Harray[53][248], Harray[54][248], Harray[55][248], Harray[56][248], Harray[57][248], Harray[58][248], Harray[59][248], Harray[60][248], Harray[61][248], Harray[62][248], Harray[63][248], Harray[64][248], Harray[65][248], Harray[66][248], Harray[67][248], Harray[68][248], Harray[69][248], Harray[70][248], Harray[71][248], Harray[72][248], Harray[73][248], Harray[74][248], Harray[75][248], Harray[76][248], Harray[77][248], Harray[78][248], Harray[79][248], Harray[80][248], Harray[81][248], Harray[82][248], Harray[83][248], Harray[84][248], Harray[85][248], Harray[86][248], Harray[87][248], Harray[88][248], Harray[89][248], Harray[90][248], Harray[91][248], Harray[92][248], Harray[93][248], Harray[94][248], Harray[95][248], Harray[96][248], Harray[97][248], Harray[98][248], Harray[99][248], Harray[100][248], Harray[101][248], Harray[102][248], Harray[103][248], Harray[104][248], Harray[105][248], Harray[106][248], Harray[107][248], Harray[108][248], Harray[109][248], Harray[110][248], Harray[111][248], Harray[112][248], Harray[113][248], Harray[114][248], Harray[115][248], Harray[116][248], Harray[117][248], Harray[118][248], Harray[119][248], Harray[120][248], Harray[121][248], Harray[122][248], Harray[123][248], Harray[124][248], Harray[125][248], Harray[126][248], Harray[127][248]};
assign h_col_249 = {Harray[0][249], Harray[1][249], Harray[2][249], Harray[3][249], Harray[4][249], Harray[5][249], Harray[6][249], Harray[7][249], Harray[8][249], Harray[9][249], Harray[10][249], Harray[11][249], Harray[12][249], Harray[13][249], Harray[14][249], Harray[15][249], Harray[16][249], Harray[17][249], Harray[18][249], Harray[19][249], Harray[20][249], Harray[21][249], Harray[22][249], Harray[23][249], Harray[24][249], Harray[25][249], Harray[26][249], Harray[27][249], Harray[28][249], Harray[29][249], Harray[30][249], Harray[31][249], Harray[32][249], Harray[33][249], Harray[34][249], Harray[35][249], Harray[36][249], Harray[37][249], Harray[38][249], Harray[39][249], Harray[40][249], Harray[41][249], Harray[42][249], Harray[43][249], Harray[44][249], Harray[45][249], Harray[46][249], Harray[47][249], Harray[48][249], Harray[49][249], Harray[50][249], Harray[51][249], Harray[52][249], Harray[53][249], Harray[54][249], Harray[55][249], Harray[56][249], Harray[57][249], Harray[58][249], Harray[59][249], Harray[60][249], Harray[61][249], Harray[62][249], Harray[63][249], Harray[64][249], Harray[65][249], Harray[66][249], Harray[67][249], Harray[68][249], Harray[69][249], Harray[70][249], Harray[71][249], Harray[72][249], Harray[73][249], Harray[74][249], Harray[75][249], Harray[76][249], Harray[77][249], Harray[78][249], Harray[79][249], Harray[80][249], Harray[81][249], Harray[82][249], Harray[83][249], Harray[84][249], Harray[85][249], Harray[86][249], Harray[87][249], Harray[88][249], Harray[89][249], Harray[90][249], Harray[91][249], Harray[92][249], Harray[93][249], Harray[94][249], Harray[95][249], Harray[96][249], Harray[97][249], Harray[98][249], Harray[99][249], Harray[100][249], Harray[101][249], Harray[102][249], Harray[103][249], Harray[104][249], Harray[105][249], Harray[106][249], Harray[107][249], Harray[108][249], Harray[109][249], Harray[110][249], Harray[111][249], Harray[112][249], Harray[113][249], Harray[114][249], Harray[115][249], Harray[116][249], Harray[117][249], Harray[118][249], Harray[119][249], Harray[120][249], Harray[121][249], Harray[122][249], Harray[123][249], Harray[124][249], Harray[125][249], Harray[126][249], Harray[127][249]};
assign h_col_250 = {Harray[0][250], Harray[1][250], Harray[2][250], Harray[3][250], Harray[4][250], Harray[5][250], Harray[6][250], Harray[7][250], Harray[8][250], Harray[9][250], Harray[10][250], Harray[11][250], Harray[12][250], Harray[13][250], Harray[14][250], Harray[15][250], Harray[16][250], Harray[17][250], Harray[18][250], Harray[19][250], Harray[20][250], Harray[21][250], Harray[22][250], Harray[23][250], Harray[24][250], Harray[25][250], Harray[26][250], Harray[27][250], Harray[28][250], Harray[29][250], Harray[30][250], Harray[31][250], Harray[32][250], Harray[33][250], Harray[34][250], Harray[35][250], Harray[36][250], Harray[37][250], Harray[38][250], Harray[39][250], Harray[40][250], Harray[41][250], Harray[42][250], Harray[43][250], Harray[44][250], Harray[45][250], Harray[46][250], Harray[47][250], Harray[48][250], Harray[49][250], Harray[50][250], Harray[51][250], Harray[52][250], Harray[53][250], Harray[54][250], Harray[55][250], Harray[56][250], Harray[57][250], Harray[58][250], Harray[59][250], Harray[60][250], Harray[61][250], Harray[62][250], Harray[63][250], Harray[64][250], Harray[65][250], Harray[66][250], Harray[67][250], Harray[68][250], Harray[69][250], Harray[70][250], Harray[71][250], Harray[72][250], Harray[73][250], Harray[74][250], Harray[75][250], Harray[76][250], Harray[77][250], Harray[78][250], Harray[79][250], Harray[80][250], Harray[81][250], Harray[82][250], Harray[83][250], Harray[84][250], Harray[85][250], Harray[86][250], Harray[87][250], Harray[88][250], Harray[89][250], Harray[90][250], Harray[91][250], Harray[92][250], Harray[93][250], Harray[94][250], Harray[95][250], Harray[96][250], Harray[97][250], Harray[98][250], Harray[99][250], Harray[100][250], Harray[101][250], Harray[102][250], Harray[103][250], Harray[104][250], Harray[105][250], Harray[106][250], Harray[107][250], Harray[108][250], Harray[109][250], Harray[110][250], Harray[111][250], Harray[112][250], Harray[113][250], Harray[114][250], Harray[115][250], Harray[116][250], Harray[117][250], Harray[118][250], Harray[119][250], Harray[120][250], Harray[121][250], Harray[122][250], Harray[123][250], Harray[124][250], Harray[125][250], Harray[126][250], Harray[127][250]};
assign h_col_251 = {Harray[0][251], Harray[1][251], Harray[2][251], Harray[3][251], Harray[4][251], Harray[5][251], Harray[6][251], Harray[7][251], Harray[8][251], Harray[9][251], Harray[10][251], Harray[11][251], Harray[12][251], Harray[13][251], Harray[14][251], Harray[15][251], Harray[16][251], Harray[17][251], Harray[18][251], Harray[19][251], Harray[20][251], Harray[21][251], Harray[22][251], Harray[23][251], Harray[24][251], Harray[25][251], Harray[26][251], Harray[27][251], Harray[28][251], Harray[29][251], Harray[30][251], Harray[31][251], Harray[32][251], Harray[33][251], Harray[34][251], Harray[35][251], Harray[36][251], Harray[37][251], Harray[38][251], Harray[39][251], Harray[40][251], Harray[41][251], Harray[42][251], Harray[43][251], Harray[44][251], Harray[45][251], Harray[46][251], Harray[47][251], Harray[48][251], Harray[49][251], Harray[50][251], Harray[51][251], Harray[52][251], Harray[53][251], Harray[54][251], Harray[55][251], Harray[56][251], Harray[57][251], Harray[58][251], Harray[59][251], Harray[60][251], Harray[61][251], Harray[62][251], Harray[63][251], Harray[64][251], Harray[65][251], Harray[66][251], Harray[67][251], Harray[68][251], Harray[69][251], Harray[70][251], Harray[71][251], Harray[72][251], Harray[73][251], Harray[74][251], Harray[75][251], Harray[76][251], Harray[77][251], Harray[78][251], Harray[79][251], Harray[80][251], Harray[81][251], Harray[82][251], Harray[83][251], Harray[84][251], Harray[85][251], Harray[86][251], Harray[87][251], Harray[88][251], Harray[89][251], Harray[90][251], Harray[91][251], Harray[92][251], Harray[93][251], Harray[94][251], Harray[95][251], Harray[96][251], Harray[97][251], Harray[98][251], Harray[99][251], Harray[100][251], Harray[101][251], Harray[102][251], Harray[103][251], Harray[104][251], Harray[105][251], Harray[106][251], Harray[107][251], Harray[108][251], Harray[109][251], Harray[110][251], Harray[111][251], Harray[112][251], Harray[113][251], Harray[114][251], Harray[115][251], Harray[116][251], Harray[117][251], Harray[118][251], Harray[119][251], Harray[120][251], Harray[121][251], Harray[122][251], Harray[123][251], Harray[124][251], Harray[125][251], Harray[126][251], Harray[127][251]};
assign h_col_252 = {Harray[0][252], Harray[1][252], Harray[2][252], Harray[3][252], Harray[4][252], Harray[5][252], Harray[6][252], Harray[7][252], Harray[8][252], Harray[9][252], Harray[10][252], Harray[11][252], Harray[12][252], Harray[13][252], Harray[14][252], Harray[15][252], Harray[16][252], Harray[17][252], Harray[18][252], Harray[19][252], Harray[20][252], Harray[21][252], Harray[22][252], Harray[23][252], Harray[24][252], Harray[25][252], Harray[26][252], Harray[27][252], Harray[28][252], Harray[29][252], Harray[30][252], Harray[31][252], Harray[32][252], Harray[33][252], Harray[34][252], Harray[35][252], Harray[36][252], Harray[37][252], Harray[38][252], Harray[39][252], Harray[40][252], Harray[41][252], Harray[42][252], Harray[43][252], Harray[44][252], Harray[45][252], Harray[46][252], Harray[47][252], Harray[48][252], Harray[49][252], Harray[50][252], Harray[51][252], Harray[52][252], Harray[53][252], Harray[54][252], Harray[55][252], Harray[56][252], Harray[57][252], Harray[58][252], Harray[59][252], Harray[60][252], Harray[61][252], Harray[62][252], Harray[63][252], Harray[64][252], Harray[65][252], Harray[66][252], Harray[67][252], Harray[68][252], Harray[69][252], Harray[70][252], Harray[71][252], Harray[72][252], Harray[73][252], Harray[74][252], Harray[75][252], Harray[76][252], Harray[77][252], Harray[78][252], Harray[79][252], Harray[80][252], Harray[81][252], Harray[82][252], Harray[83][252], Harray[84][252], Harray[85][252], Harray[86][252], Harray[87][252], Harray[88][252], Harray[89][252], Harray[90][252], Harray[91][252], Harray[92][252], Harray[93][252], Harray[94][252], Harray[95][252], Harray[96][252], Harray[97][252], Harray[98][252], Harray[99][252], Harray[100][252], Harray[101][252], Harray[102][252], Harray[103][252], Harray[104][252], Harray[105][252], Harray[106][252], Harray[107][252], Harray[108][252], Harray[109][252], Harray[110][252], Harray[111][252], Harray[112][252], Harray[113][252], Harray[114][252], Harray[115][252], Harray[116][252], Harray[117][252], Harray[118][252], Harray[119][252], Harray[120][252], Harray[121][252], Harray[122][252], Harray[123][252], Harray[124][252], Harray[125][252], Harray[126][252], Harray[127][252]};
assign h_col_253 = {Harray[0][253], Harray[1][253], Harray[2][253], Harray[3][253], Harray[4][253], Harray[5][253], Harray[6][253], Harray[7][253], Harray[8][253], Harray[9][253], Harray[10][253], Harray[11][253], Harray[12][253], Harray[13][253], Harray[14][253], Harray[15][253], Harray[16][253], Harray[17][253], Harray[18][253], Harray[19][253], Harray[20][253], Harray[21][253], Harray[22][253], Harray[23][253], Harray[24][253], Harray[25][253], Harray[26][253], Harray[27][253], Harray[28][253], Harray[29][253], Harray[30][253], Harray[31][253], Harray[32][253], Harray[33][253], Harray[34][253], Harray[35][253], Harray[36][253], Harray[37][253], Harray[38][253], Harray[39][253], Harray[40][253], Harray[41][253], Harray[42][253], Harray[43][253], Harray[44][253], Harray[45][253], Harray[46][253], Harray[47][253], Harray[48][253], Harray[49][253], Harray[50][253], Harray[51][253], Harray[52][253], Harray[53][253], Harray[54][253], Harray[55][253], Harray[56][253], Harray[57][253], Harray[58][253], Harray[59][253], Harray[60][253], Harray[61][253], Harray[62][253], Harray[63][253], Harray[64][253], Harray[65][253], Harray[66][253], Harray[67][253], Harray[68][253], Harray[69][253], Harray[70][253], Harray[71][253], Harray[72][253], Harray[73][253], Harray[74][253], Harray[75][253], Harray[76][253], Harray[77][253], Harray[78][253], Harray[79][253], Harray[80][253], Harray[81][253], Harray[82][253], Harray[83][253], Harray[84][253], Harray[85][253], Harray[86][253], Harray[87][253], Harray[88][253], Harray[89][253], Harray[90][253], Harray[91][253], Harray[92][253], Harray[93][253], Harray[94][253], Harray[95][253], Harray[96][253], Harray[97][253], Harray[98][253], Harray[99][253], Harray[100][253], Harray[101][253], Harray[102][253], Harray[103][253], Harray[104][253], Harray[105][253], Harray[106][253], Harray[107][253], Harray[108][253], Harray[109][253], Harray[110][253], Harray[111][253], Harray[112][253], Harray[113][253], Harray[114][253], Harray[115][253], Harray[116][253], Harray[117][253], Harray[118][253], Harray[119][253], Harray[120][253], Harray[121][253], Harray[122][253], Harray[123][253], Harray[124][253], Harray[125][253], Harray[126][253], Harray[127][253]};
assign h_col_254 = {Harray[0][254], Harray[1][254], Harray[2][254], Harray[3][254], Harray[4][254], Harray[5][254], Harray[6][254], Harray[7][254], Harray[8][254], Harray[9][254], Harray[10][254], Harray[11][254], Harray[12][254], Harray[13][254], Harray[14][254], Harray[15][254], Harray[16][254], Harray[17][254], Harray[18][254], Harray[19][254], Harray[20][254], Harray[21][254], Harray[22][254], Harray[23][254], Harray[24][254], Harray[25][254], Harray[26][254], Harray[27][254], Harray[28][254], Harray[29][254], Harray[30][254], Harray[31][254], Harray[32][254], Harray[33][254], Harray[34][254], Harray[35][254], Harray[36][254], Harray[37][254], Harray[38][254], Harray[39][254], Harray[40][254], Harray[41][254], Harray[42][254], Harray[43][254], Harray[44][254], Harray[45][254], Harray[46][254], Harray[47][254], Harray[48][254], Harray[49][254], Harray[50][254], Harray[51][254], Harray[52][254], Harray[53][254], Harray[54][254], Harray[55][254], Harray[56][254], Harray[57][254], Harray[58][254], Harray[59][254], Harray[60][254], Harray[61][254], Harray[62][254], Harray[63][254], Harray[64][254], Harray[65][254], Harray[66][254], Harray[67][254], Harray[68][254], Harray[69][254], Harray[70][254], Harray[71][254], Harray[72][254], Harray[73][254], Harray[74][254], Harray[75][254], Harray[76][254], Harray[77][254], Harray[78][254], Harray[79][254], Harray[80][254], Harray[81][254], Harray[82][254], Harray[83][254], Harray[84][254], Harray[85][254], Harray[86][254], Harray[87][254], Harray[88][254], Harray[89][254], Harray[90][254], Harray[91][254], Harray[92][254], Harray[93][254], Harray[94][254], Harray[95][254], Harray[96][254], Harray[97][254], Harray[98][254], Harray[99][254], Harray[100][254], Harray[101][254], Harray[102][254], Harray[103][254], Harray[104][254], Harray[105][254], Harray[106][254], Harray[107][254], Harray[108][254], Harray[109][254], Harray[110][254], Harray[111][254], Harray[112][254], Harray[113][254], Harray[114][254], Harray[115][254], Harray[116][254], Harray[117][254], Harray[118][254], Harray[119][254], Harray[120][254], Harray[121][254], Harray[122][254], Harray[123][254], Harray[124][254], Harray[125][254], Harray[126][254], Harray[127][254]};
assign h_col_255 = {Harray[0][255], Harray[1][255], Harray[2][255], Harray[3][255], Harray[4][255], Harray[5][255], Harray[6][255], Harray[7][255], Harray[8][255], Harray[9][255], Harray[10][255], Harray[11][255], Harray[12][255], Harray[13][255], Harray[14][255], Harray[15][255], Harray[16][255], Harray[17][255], Harray[18][255], Harray[19][255], Harray[20][255], Harray[21][255], Harray[22][255], Harray[23][255], Harray[24][255], Harray[25][255], Harray[26][255], Harray[27][255], Harray[28][255], Harray[29][255], Harray[30][255], Harray[31][255], Harray[32][255], Harray[33][255], Harray[34][255], Harray[35][255], Harray[36][255], Harray[37][255], Harray[38][255], Harray[39][255], Harray[40][255], Harray[41][255], Harray[42][255], Harray[43][255], Harray[44][255], Harray[45][255], Harray[46][255], Harray[47][255], Harray[48][255], Harray[49][255], Harray[50][255], Harray[51][255], Harray[52][255], Harray[53][255], Harray[54][255], Harray[55][255], Harray[56][255], Harray[57][255], Harray[58][255], Harray[59][255], Harray[60][255], Harray[61][255], Harray[62][255], Harray[63][255], Harray[64][255], Harray[65][255], Harray[66][255], Harray[67][255], Harray[68][255], Harray[69][255], Harray[70][255], Harray[71][255], Harray[72][255], Harray[73][255], Harray[74][255], Harray[75][255], Harray[76][255], Harray[77][255], Harray[78][255], Harray[79][255], Harray[80][255], Harray[81][255], Harray[82][255], Harray[83][255], Harray[84][255], Harray[85][255], Harray[86][255], Harray[87][255], Harray[88][255], Harray[89][255], Harray[90][255], Harray[91][255], Harray[92][255], Harray[93][255], Harray[94][255], Harray[95][255], Harray[96][255], Harray[97][255], Harray[98][255], Harray[99][255], Harray[100][255], Harray[101][255], Harray[102][255], Harray[103][255], Harray[104][255], Harray[105][255], Harray[106][255], Harray[107][255], Harray[108][255], Harray[109][255], Harray[110][255], Harray[111][255], Harray[112][255], Harray[113][255], Harray[114][255], Harray[115][255], Harray[116][255], Harray[117][255], Harray[118][255], Harray[119][255], Harray[120][255], Harray[121][255], Harray[122][255], Harray[123][255], Harray[124][255], Harray[125][255], Harray[126][255], Harray[127][255]};


wire [7:0] check_col_0, check_col_1, check_col_2, check_col_3, check_col_4, check_col_5, check_col_6, check_col_7, 
           check_col_8, check_col_9, check_col_10, check_col_11, check_col_12, check_col_13, check_col_14, check_col_15, 
           check_col_16, check_col_17, check_col_18, check_col_19, check_col_20, check_col_21, check_col_22, check_col_23, 
           check_col_24, check_col_25, check_col_26, check_col_27, check_col_28, check_col_29, check_col_30, check_col_31, 
           check_col_32, check_col_33, check_col_34, check_col_35, check_col_36, check_col_37, check_col_38, check_col_39, 
           check_col_40, check_col_41, check_col_42, check_col_43, check_col_44, check_col_45, check_col_46, check_col_47, 
           check_col_48, check_col_49, check_col_50, check_col_51, check_col_52, check_col_53, check_col_54, check_col_55, 
           check_col_56, check_col_57, check_col_58, check_col_59, check_col_60, check_col_61, check_col_62, check_col_63, 
           check_col_64, check_col_65, check_col_66, check_col_67, check_col_68, check_col_69, check_col_70, check_col_71, 
           check_col_72, check_col_73, check_col_74, check_col_75, check_col_76, check_col_77, check_col_78, check_col_79, 
           check_col_80, check_col_81, check_col_82, check_col_83, check_col_84, check_col_85, check_col_86, check_col_87, 
           check_col_88, check_col_89, check_col_90, check_col_91, check_col_92, check_col_93, check_col_94, check_col_95, 
           check_col_96, check_col_97, check_col_98, check_col_99, check_col_100, check_col_101, check_col_102, check_col_103, 
           check_col_104, check_col_105, check_col_106, check_col_107, check_col_108, check_col_109, check_col_110, check_col_111, 
           check_col_112, check_col_113, check_col_114, check_col_115, check_col_116, check_col_117, check_col_118, check_col_119, 
           check_col_120, check_col_121, check_col_122, check_col_123, check_col_124, check_col_125, check_col_126, check_col_127, 
           check_col_128, check_col_129, check_col_130, check_col_131, check_col_132, check_col_133, check_col_134, check_col_135, 
           check_col_136, check_col_137, check_col_138, check_col_139, check_col_140, check_col_141, check_col_142, check_col_143, 
           check_col_144, check_col_145, check_col_146, check_col_147, check_col_148, check_col_149, check_col_150, check_col_151, 
           check_col_152, check_col_153, check_col_154, check_col_155, check_col_156, check_col_157, check_col_158, check_col_159, 
           check_col_160, check_col_161, check_col_162, check_col_163, check_col_164, check_col_165, check_col_166, check_col_167, 
           check_col_168, check_col_169, check_col_170, check_col_171, check_col_172, check_col_173, check_col_174, check_col_175, 
           check_col_176, check_col_177, check_col_178, check_col_179, check_col_180, check_col_181, check_col_182, check_col_183, 
           check_col_184, check_col_185, check_col_186, check_col_187, check_col_188, check_col_189, check_col_190, check_col_191, 
           check_col_192, check_col_193, check_col_194, check_col_195, check_col_196, check_col_197, check_col_198, check_col_199, 
           check_col_200, check_col_201, check_col_202, check_col_203, check_col_204, check_col_205, check_col_206, check_col_207, 
           check_col_208, check_col_209, check_col_210, check_col_211, check_col_212, check_col_213, check_col_214, check_col_215, 
           check_col_216, check_col_217, check_col_218, check_col_219, check_col_220, check_col_221, check_col_222, check_col_223, 
           check_col_224, check_col_225, check_col_226, check_col_227, check_col_228, check_col_229, check_col_230, check_col_231, 
           check_col_232, check_col_233, check_col_234, check_col_235, check_col_236, check_col_237, check_col_238, check_col_239, 
           check_col_240, check_col_241, check_col_242, check_col_243, check_col_244, check_col_245, check_col_246, check_col_247, 
           check_col_248, check_col_249, check_col_250, check_col_251, check_col_252, check_col_253, check_col_254, check_col_255;

wire [7:0] wrong_col_0, wrong_col_1, wrong_col_2, wrong_col_3, wrong_col_4, wrong_col_5, wrong_col_6, wrong_col_7, 
           wrong_col_8, wrong_col_9, wrong_col_10, wrong_col_11, wrong_col_12, wrong_col_13, wrong_col_14, wrong_col_15, 
           wrong_col_16, wrong_col_17, wrong_col_18, wrong_col_19, wrong_col_20, wrong_col_21, wrong_col_22, wrong_col_23, 
           wrong_col_24, wrong_col_25, wrong_col_26, wrong_col_27, wrong_col_28, wrong_col_29, wrong_col_30, wrong_col_31, 
           wrong_col_32, wrong_col_33, wrong_col_34, wrong_col_35, wrong_col_36, wrong_col_37, wrong_col_38, wrong_col_39, 
           wrong_col_40, wrong_col_41, wrong_col_42, wrong_col_43, wrong_col_44, wrong_col_45, wrong_col_46, wrong_col_47, 
           wrong_col_48, wrong_col_49, wrong_col_50, wrong_col_51, wrong_col_52, wrong_col_53, wrong_col_54, wrong_col_55, 
           wrong_col_56, wrong_col_57, wrong_col_58, wrong_col_59, wrong_col_60, wrong_col_61, wrong_col_62, wrong_col_63, 
           wrong_col_64, wrong_col_65, wrong_col_66, wrong_col_67, wrong_col_68, wrong_col_69, wrong_col_70, wrong_col_71, 
           wrong_col_72, wrong_col_73, wrong_col_74, wrong_col_75, wrong_col_76, wrong_col_77, wrong_col_78, wrong_col_79, 
           wrong_col_80, wrong_col_81, wrong_col_82, wrong_col_83, wrong_col_84, wrong_col_85, wrong_col_86, wrong_col_87, 
           wrong_col_88, wrong_col_89, wrong_col_90, wrong_col_91, wrong_col_92, wrong_col_93, wrong_col_94, wrong_col_95, 
           wrong_col_96, wrong_col_97, wrong_col_98, wrong_col_99, wrong_col_100, wrong_col_101, wrong_col_102, wrong_col_103, 
           wrong_col_104, wrong_col_105, wrong_col_106, wrong_col_107, wrong_col_108, wrong_col_109, wrong_col_110, wrong_col_111, 
           wrong_col_112, wrong_col_113, wrong_col_114, wrong_col_115, wrong_col_116, wrong_col_117, wrong_col_118, wrong_col_119, 
           wrong_col_120, wrong_col_121, wrong_col_122, wrong_col_123, wrong_col_124, wrong_col_125, wrong_col_126, wrong_col_127, 
           wrong_col_128, wrong_col_129, wrong_col_130, wrong_col_131, wrong_col_132, wrong_col_133, wrong_col_134, wrong_col_135, 
           wrong_col_136, wrong_col_137, wrong_col_138, wrong_col_139, wrong_col_140, wrong_col_141, wrong_col_142, wrong_col_143, 
           wrong_col_144, wrong_col_145, wrong_col_146, wrong_col_147, wrong_col_148, wrong_col_149, wrong_col_150, wrong_col_151, 
           wrong_col_152, wrong_col_153, wrong_col_154, wrong_col_155, wrong_col_156, wrong_col_157, wrong_col_158, wrong_col_159, 
           wrong_col_160, wrong_col_161, wrong_col_162, wrong_col_163, wrong_col_164, wrong_col_165, wrong_col_166, wrong_col_167, 
           wrong_col_168, wrong_col_169, wrong_col_170, wrong_col_171, wrong_col_172, wrong_col_173, wrong_col_174, wrong_col_175, 
           wrong_col_176, wrong_col_177, wrong_col_178, wrong_col_179, wrong_col_180, wrong_col_181, wrong_col_182, wrong_col_183, 
           wrong_col_184, wrong_col_185, wrong_col_186, wrong_col_187, wrong_col_188, wrong_col_189, wrong_col_190, wrong_col_191, 
           wrong_col_192, wrong_col_193, wrong_col_194, wrong_col_195, wrong_col_196, wrong_col_197, wrong_col_198, wrong_col_199, 
           wrong_col_200, wrong_col_201, wrong_col_202, wrong_col_203, wrong_col_204, wrong_col_205, wrong_col_206, wrong_col_207, 
           wrong_col_208, wrong_col_209, wrong_col_210, wrong_col_211, wrong_col_212, wrong_col_213, wrong_col_214, wrong_col_215, 
           wrong_col_216, wrong_col_217, wrong_col_218, wrong_col_219, wrong_col_220, wrong_col_221, wrong_col_222, wrong_col_223, 
           wrong_col_224, wrong_col_225, wrong_col_226, wrong_col_227, wrong_col_228, wrong_col_229, wrong_col_230, wrong_col_231, 
           wrong_col_232, wrong_col_233, wrong_col_234, wrong_col_235, wrong_col_236, wrong_col_237, wrong_col_238, wrong_col_239, 
           wrong_col_240, wrong_col_241, wrong_col_242, wrong_col_243, wrong_col_244, wrong_col_245, wrong_col_246, wrong_col_247, 
           wrong_col_248, wrong_col_249, wrong_col_250, wrong_col_251, wrong_col_252, wrong_col_253, wrong_col_254, wrong_col_255;

bitsadder_128 c_num_0(.data_in(h_col_0), .sum(check_col_0));
bitsadder_128 c_num_1(.data_in(h_col_1), .sum(check_col_1));
bitsadder_128 c_num_2(.data_in(h_col_2), .sum(check_col_2));
bitsadder_128 c_num_3(.data_in(h_col_3), .sum(check_col_3));
bitsadder_128 c_num_4(.data_in(h_col_4), .sum(check_col_4));
bitsadder_128 c_num_5(.data_in(h_col_5), .sum(check_col_5));
bitsadder_128 c_num_6(.data_in(h_col_6), .sum(check_col_6));
bitsadder_128 c_num_7(.data_in(h_col_7), .sum(check_col_7));
bitsadder_128 c_num_8(.data_in(h_col_8), .sum(check_col_8));
bitsadder_128 c_num_9(.data_in(h_col_9), .sum(check_col_9));
bitsadder_128 c_num_10(.data_in(h_col_10), .sum(check_col_10));
bitsadder_128 c_num_11(.data_in(h_col_11), .sum(check_col_11));
bitsadder_128 c_num_12(.data_in(h_col_12), .sum(check_col_12));
bitsadder_128 c_num_13(.data_in(h_col_13), .sum(check_col_13));
bitsadder_128 c_num_14(.data_in(h_col_14), .sum(check_col_14));
bitsadder_128 c_num_15(.data_in(h_col_15), .sum(check_col_15));
bitsadder_128 c_num_16(.data_in(h_col_16), .sum(check_col_16));
bitsadder_128 c_num_17(.data_in(h_col_17), .sum(check_col_17));
bitsadder_128 c_num_18(.data_in(h_col_18), .sum(check_col_18));
bitsadder_128 c_num_19(.data_in(h_col_19), .sum(check_col_19));
bitsadder_128 c_num_20(.data_in(h_col_20), .sum(check_col_20));
bitsadder_128 c_num_21(.data_in(h_col_21), .sum(check_col_21));
bitsadder_128 c_num_22(.data_in(h_col_22), .sum(check_col_22));
bitsadder_128 c_num_23(.data_in(h_col_23), .sum(check_col_23));
bitsadder_128 c_num_24(.data_in(h_col_24), .sum(check_col_24));
bitsadder_128 c_num_25(.data_in(h_col_25), .sum(check_col_25));
bitsadder_128 c_num_26(.data_in(h_col_26), .sum(check_col_26));
bitsadder_128 c_num_27(.data_in(h_col_27), .sum(check_col_27));
bitsadder_128 c_num_28(.data_in(h_col_28), .sum(check_col_28));
bitsadder_128 c_num_29(.data_in(h_col_29), .sum(check_col_29));
bitsadder_128 c_num_30(.data_in(h_col_30), .sum(check_col_30));
bitsadder_128 c_num_31(.data_in(h_col_31), .sum(check_col_31));
bitsadder_128 c_num_32(.data_in(h_col_32), .sum(check_col_32));
bitsadder_128 c_num_33(.data_in(h_col_33), .sum(check_col_33));
bitsadder_128 c_num_34(.data_in(h_col_34), .sum(check_col_34));
bitsadder_128 c_num_35(.data_in(h_col_35), .sum(check_col_35));
bitsadder_128 c_num_36(.data_in(h_col_36), .sum(check_col_36));
bitsadder_128 c_num_37(.data_in(h_col_37), .sum(check_col_37));
bitsadder_128 c_num_38(.data_in(h_col_38), .sum(check_col_38));
bitsadder_128 c_num_39(.data_in(h_col_39), .sum(check_col_39));
bitsadder_128 c_num_40(.data_in(h_col_40), .sum(check_col_40));
bitsadder_128 c_num_41(.data_in(h_col_41), .sum(check_col_41));
bitsadder_128 c_num_42(.data_in(h_col_42), .sum(check_col_42));
bitsadder_128 c_num_43(.data_in(h_col_43), .sum(check_col_43));
bitsadder_128 c_num_44(.data_in(h_col_44), .sum(check_col_44));
bitsadder_128 c_num_45(.data_in(h_col_45), .sum(check_col_45));
bitsadder_128 c_num_46(.data_in(h_col_46), .sum(check_col_46));
bitsadder_128 c_num_47(.data_in(h_col_47), .sum(check_col_47));
bitsadder_128 c_num_48(.data_in(h_col_48), .sum(check_col_48));
bitsadder_128 c_num_49(.data_in(h_col_49), .sum(check_col_49));
bitsadder_128 c_num_50(.data_in(h_col_50), .sum(check_col_50));
bitsadder_128 c_num_51(.data_in(h_col_51), .sum(check_col_51));
bitsadder_128 c_num_52(.data_in(h_col_52), .sum(check_col_52));
bitsadder_128 c_num_53(.data_in(h_col_53), .sum(check_col_53));
bitsadder_128 c_num_54(.data_in(h_col_54), .sum(check_col_54));
bitsadder_128 c_num_55(.data_in(h_col_55), .sum(check_col_55));
bitsadder_128 c_num_56(.data_in(h_col_56), .sum(check_col_56));
bitsadder_128 c_num_57(.data_in(h_col_57), .sum(check_col_57));
bitsadder_128 c_num_58(.data_in(h_col_58), .sum(check_col_58));
bitsadder_128 c_num_59(.data_in(h_col_59), .sum(check_col_59));
bitsadder_128 c_num_60(.data_in(h_col_60), .sum(check_col_60));
bitsadder_128 c_num_61(.data_in(h_col_61), .sum(check_col_61));
bitsadder_128 c_num_62(.data_in(h_col_62), .sum(check_col_62));
bitsadder_128 c_num_63(.data_in(h_col_63), .sum(check_col_63));
bitsadder_128 c_num_64(.data_in(h_col_64), .sum(check_col_64));
bitsadder_128 c_num_65(.data_in(h_col_65), .sum(check_col_65));
bitsadder_128 c_num_66(.data_in(h_col_66), .sum(check_col_66));
bitsadder_128 c_num_67(.data_in(h_col_67), .sum(check_col_67));
bitsadder_128 c_num_68(.data_in(h_col_68), .sum(check_col_68));
bitsadder_128 c_num_69(.data_in(h_col_69), .sum(check_col_69));
bitsadder_128 c_num_70(.data_in(h_col_70), .sum(check_col_70));
bitsadder_128 c_num_71(.data_in(h_col_71), .sum(check_col_71));
bitsadder_128 c_num_72(.data_in(h_col_72), .sum(check_col_72));
bitsadder_128 c_num_73(.data_in(h_col_73), .sum(check_col_73));
bitsadder_128 c_num_74(.data_in(h_col_74), .sum(check_col_74));
bitsadder_128 c_num_75(.data_in(h_col_75), .sum(check_col_75));
bitsadder_128 c_num_76(.data_in(h_col_76), .sum(check_col_76));
bitsadder_128 c_num_77(.data_in(h_col_77), .sum(check_col_77));
bitsadder_128 c_num_78(.data_in(h_col_78), .sum(check_col_78));
bitsadder_128 c_num_79(.data_in(h_col_79), .sum(check_col_79));
bitsadder_128 c_num_80(.data_in(h_col_80), .sum(check_col_80));
bitsadder_128 c_num_81(.data_in(h_col_81), .sum(check_col_81));
bitsadder_128 c_num_82(.data_in(h_col_82), .sum(check_col_82));
bitsadder_128 c_num_83(.data_in(h_col_83), .sum(check_col_83));
bitsadder_128 c_num_84(.data_in(h_col_84), .sum(check_col_84));
bitsadder_128 c_num_85(.data_in(h_col_85), .sum(check_col_85));
bitsadder_128 c_num_86(.data_in(h_col_86), .sum(check_col_86));
bitsadder_128 c_num_87(.data_in(h_col_87), .sum(check_col_87));
bitsadder_128 c_num_88(.data_in(h_col_88), .sum(check_col_88));
bitsadder_128 c_num_89(.data_in(h_col_89), .sum(check_col_89));
bitsadder_128 c_num_90(.data_in(h_col_90), .sum(check_col_90));
bitsadder_128 c_num_91(.data_in(h_col_91), .sum(check_col_91));
bitsadder_128 c_num_92(.data_in(h_col_92), .sum(check_col_92));
bitsadder_128 c_num_93(.data_in(h_col_93), .sum(check_col_93));
bitsadder_128 c_num_94(.data_in(h_col_94), .sum(check_col_94));
bitsadder_128 c_num_95(.data_in(h_col_95), .sum(check_col_95));
bitsadder_128 c_num_96(.data_in(h_col_96), .sum(check_col_96));
bitsadder_128 c_num_97(.data_in(h_col_97), .sum(check_col_97));
bitsadder_128 c_num_98(.data_in(h_col_98), .sum(check_col_98));
bitsadder_128 c_num_99(.data_in(h_col_99), .sum(check_col_99));
bitsadder_128 c_num_100(.data_in(h_col_100), .sum(check_col_100));
bitsadder_128 c_num_101(.data_in(h_col_101), .sum(check_col_101));
bitsadder_128 c_num_102(.data_in(h_col_102), .sum(check_col_102));
bitsadder_128 c_num_103(.data_in(h_col_103), .sum(check_col_103));
bitsadder_128 c_num_104(.data_in(h_col_104), .sum(check_col_104));
bitsadder_128 c_num_105(.data_in(h_col_105), .sum(check_col_105));
bitsadder_128 c_num_106(.data_in(h_col_106), .sum(check_col_106));
bitsadder_128 c_num_107(.data_in(h_col_107), .sum(check_col_107));
bitsadder_128 c_num_108(.data_in(h_col_108), .sum(check_col_108));
bitsadder_128 c_num_109(.data_in(h_col_109), .sum(check_col_109));
bitsadder_128 c_num_110(.data_in(h_col_110), .sum(check_col_110));
bitsadder_128 c_num_111(.data_in(h_col_111), .sum(check_col_111));
bitsadder_128 c_num_112(.data_in(h_col_112), .sum(check_col_112));
bitsadder_128 c_num_113(.data_in(h_col_113), .sum(check_col_113));
bitsadder_128 c_num_114(.data_in(h_col_114), .sum(check_col_114));
bitsadder_128 c_num_115(.data_in(h_col_115), .sum(check_col_115));
bitsadder_128 c_num_116(.data_in(h_col_116), .sum(check_col_116));
bitsadder_128 c_num_117(.data_in(h_col_117), .sum(check_col_117));
bitsadder_128 c_num_118(.data_in(h_col_118), .sum(check_col_118));
bitsadder_128 c_num_119(.data_in(h_col_119), .sum(check_col_119));
bitsadder_128 c_num_120(.data_in(h_col_120), .sum(check_col_120));
bitsadder_128 c_num_121(.data_in(h_col_121), .sum(check_col_121));
bitsadder_128 c_num_122(.data_in(h_col_122), .sum(check_col_122));
bitsadder_128 c_num_123(.data_in(h_col_123), .sum(check_col_123));
bitsadder_128 c_num_124(.data_in(h_col_124), .sum(check_col_124));
bitsadder_128 c_num_125(.data_in(h_col_125), .sum(check_col_125));
bitsadder_128 c_num_126(.data_in(h_col_126), .sum(check_col_126));
bitsadder_128 c_num_127(.data_in(h_col_127), .sum(check_col_127));
bitsadder_128 c_num_128(.data_in(h_col_128), .sum(check_col_128));
bitsadder_128 c_num_129(.data_in(h_col_129), .sum(check_col_129));
bitsadder_128 c_num_130(.data_in(h_col_130), .sum(check_col_130));
bitsadder_128 c_num_131(.data_in(h_col_131), .sum(check_col_131));
bitsadder_128 c_num_132(.data_in(h_col_132), .sum(check_col_132));
bitsadder_128 c_num_133(.data_in(h_col_133), .sum(check_col_133));
bitsadder_128 c_num_134(.data_in(h_col_134), .sum(check_col_134));
bitsadder_128 c_num_135(.data_in(h_col_135), .sum(check_col_135));
bitsadder_128 c_num_136(.data_in(h_col_136), .sum(check_col_136));
bitsadder_128 c_num_137(.data_in(h_col_137), .sum(check_col_137));
bitsadder_128 c_num_138(.data_in(h_col_138), .sum(check_col_138));
bitsadder_128 c_num_139(.data_in(h_col_139), .sum(check_col_139));
bitsadder_128 c_num_140(.data_in(h_col_140), .sum(check_col_140));
bitsadder_128 c_num_141(.data_in(h_col_141), .sum(check_col_141));
bitsadder_128 c_num_142(.data_in(h_col_142), .sum(check_col_142));
bitsadder_128 c_num_143(.data_in(h_col_143), .sum(check_col_143));
bitsadder_128 c_num_144(.data_in(h_col_144), .sum(check_col_144));
bitsadder_128 c_num_145(.data_in(h_col_145), .sum(check_col_145));
bitsadder_128 c_num_146(.data_in(h_col_146), .sum(check_col_146));
bitsadder_128 c_num_147(.data_in(h_col_147), .sum(check_col_147));
bitsadder_128 c_num_148(.data_in(h_col_148), .sum(check_col_148));
bitsadder_128 c_num_149(.data_in(h_col_149), .sum(check_col_149));
bitsadder_128 c_num_150(.data_in(h_col_150), .sum(check_col_150));
bitsadder_128 c_num_151(.data_in(h_col_151), .sum(check_col_151));
bitsadder_128 c_num_152(.data_in(h_col_152), .sum(check_col_152));
bitsadder_128 c_num_153(.data_in(h_col_153), .sum(check_col_153));
bitsadder_128 c_num_154(.data_in(h_col_154), .sum(check_col_154));
bitsadder_128 c_num_155(.data_in(h_col_155), .sum(check_col_155));
bitsadder_128 c_num_156(.data_in(h_col_156), .sum(check_col_156));
bitsadder_128 c_num_157(.data_in(h_col_157), .sum(check_col_157));
bitsadder_128 c_num_158(.data_in(h_col_158), .sum(check_col_158));
bitsadder_128 c_num_159(.data_in(h_col_159), .sum(check_col_159));
bitsadder_128 c_num_160(.data_in(h_col_160), .sum(check_col_160));
bitsadder_128 c_num_161(.data_in(h_col_161), .sum(check_col_161));
bitsadder_128 c_num_162(.data_in(h_col_162), .sum(check_col_162));
bitsadder_128 c_num_163(.data_in(h_col_163), .sum(check_col_163));
bitsadder_128 c_num_164(.data_in(h_col_164), .sum(check_col_164));
bitsadder_128 c_num_165(.data_in(h_col_165), .sum(check_col_165));
bitsadder_128 c_num_166(.data_in(h_col_166), .sum(check_col_166));
bitsadder_128 c_num_167(.data_in(h_col_167), .sum(check_col_167));
bitsadder_128 c_num_168(.data_in(h_col_168), .sum(check_col_168));
bitsadder_128 c_num_169(.data_in(h_col_169), .sum(check_col_169));
bitsadder_128 c_num_170(.data_in(h_col_170), .sum(check_col_170));
bitsadder_128 c_num_171(.data_in(h_col_171), .sum(check_col_171));
bitsadder_128 c_num_172(.data_in(h_col_172), .sum(check_col_172));
bitsadder_128 c_num_173(.data_in(h_col_173), .sum(check_col_173));
bitsadder_128 c_num_174(.data_in(h_col_174), .sum(check_col_174));
bitsadder_128 c_num_175(.data_in(h_col_175), .sum(check_col_175));
bitsadder_128 c_num_176(.data_in(h_col_176), .sum(check_col_176));
bitsadder_128 c_num_177(.data_in(h_col_177), .sum(check_col_177));
bitsadder_128 c_num_178(.data_in(h_col_178), .sum(check_col_178));
bitsadder_128 c_num_179(.data_in(h_col_179), .sum(check_col_179));
bitsadder_128 c_num_180(.data_in(h_col_180), .sum(check_col_180));
bitsadder_128 c_num_181(.data_in(h_col_181), .sum(check_col_181));
bitsadder_128 c_num_182(.data_in(h_col_182), .sum(check_col_182));
bitsadder_128 c_num_183(.data_in(h_col_183), .sum(check_col_183));
bitsadder_128 c_num_184(.data_in(h_col_184), .sum(check_col_184));
bitsadder_128 c_num_185(.data_in(h_col_185), .sum(check_col_185));
bitsadder_128 c_num_186(.data_in(h_col_186), .sum(check_col_186));
bitsadder_128 c_num_187(.data_in(h_col_187), .sum(check_col_187));
bitsadder_128 c_num_188(.data_in(h_col_188), .sum(check_col_188));
bitsadder_128 c_num_189(.data_in(h_col_189), .sum(check_col_189));
bitsadder_128 c_num_190(.data_in(h_col_190), .sum(check_col_190));
bitsadder_128 c_num_191(.data_in(h_col_191), .sum(check_col_191));
bitsadder_128 c_num_192(.data_in(h_col_192), .sum(check_col_192));
bitsadder_128 c_num_193(.data_in(h_col_193), .sum(check_col_193));
bitsadder_128 c_num_194(.data_in(h_col_194), .sum(check_col_194));
bitsadder_128 c_num_195(.data_in(h_col_195), .sum(check_col_195));
bitsadder_128 c_num_196(.data_in(h_col_196), .sum(check_col_196));
bitsadder_128 c_num_197(.data_in(h_col_197), .sum(check_col_197));
bitsadder_128 c_num_198(.data_in(h_col_198), .sum(check_col_198));
bitsadder_128 c_num_199(.data_in(h_col_199), .sum(check_col_199));
bitsadder_128 c_num_200(.data_in(h_col_200), .sum(check_col_200));
bitsadder_128 c_num_201(.data_in(h_col_201), .sum(check_col_201));
bitsadder_128 c_num_202(.data_in(h_col_202), .sum(check_col_202));
bitsadder_128 c_num_203(.data_in(h_col_203), .sum(check_col_203));
bitsadder_128 c_num_204(.data_in(h_col_204), .sum(check_col_204));
bitsadder_128 c_num_205(.data_in(h_col_205), .sum(check_col_205));
bitsadder_128 c_num_206(.data_in(h_col_206), .sum(check_col_206));
bitsadder_128 c_num_207(.data_in(h_col_207), .sum(check_col_207));
bitsadder_128 c_num_208(.data_in(h_col_208), .sum(check_col_208));
bitsadder_128 c_num_209(.data_in(h_col_209), .sum(check_col_209));
bitsadder_128 c_num_210(.data_in(h_col_210), .sum(check_col_210));
bitsadder_128 c_num_211(.data_in(h_col_211), .sum(check_col_211));
bitsadder_128 c_num_212(.data_in(h_col_212), .sum(check_col_212));
bitsadder_128 c_num_213(.data_in(h_col_213), .sum(check_col_213));
bitsadder_128 c_num_214(.data_in(h_col_214), .sum(check_col_214));
bitsadder_128 c_num_215(.data_in(h_col_215), .sum(check_col_215));
bitsadder_128 c_num_216(.data_in(h_col_216), .sum(check_col_216));
bitsadder_128 c_num_217(.data_in(h_col_217), .sum(check_col_217));
bitsadder_128 c_num_218(.data_in(h_col_218), .sum(check_col_218));
bitsadder_128 c_num_219(.data_in(h_col_219), .sum(check_col_219));
bitsadder_128 c_num_220(.data_in(h_col_220), .sum(check_col_220));
bitsadder_128 c_num_221(.data_in(h_col_221), .sum(check_col_221));
bitsadder_128 c_num_222(.data_in(h_col_222), .sum(check_col_222));
bitsadder_128 c_num_223(.data_in(h_col_223), .sum(check_col_223));
bitsadder_128 c_num_224(.data_in(h_col_224), .sum(check_col_224));
bitsadder_128 c_num_225(.data_in(h_col_225), .sum(check_col_225));
bitsadder_128 c_num_226(.data_in(h_col_226), .sum(check_col_226));
bitsadder_128 c_num_227(.data_in(h_col_227), .sum(check_col_227));
bitsadder_128 c_num_228(.data_in(h_col_228), .sum(check_col_228));
bitsadder_128 c_num_229(.data_in(h_col_229), .sum(check_col_229));
bitsadder_128 c_num_230(.data_in(h_col_230), .sum(check_col_230));
bitsadder_128 c_num_231(.data_in(h_col_231), .sum(check_col_231));
bitsadder_128 c_num_232(.data_in(h_col_232), .sum(check_col_232));
bitsadder_128 c_num_233(.data_in(h_col_233), .sum(check_col_233));
bitsadder_128 c_num_234(.data_in(h_col_234), .sum(check_col_234));
bitsadder_128 c_num_235(.data_in(h_col_235), .sum(check_col_235));
bitsadder_128 c_num_236(.data_in(h_col_236), .sum(check_col_236));
bitsadder_128 c_num_237(.data_in(h_col_237), .sum(check_col_237));
bitsadder_128 c_num_238(.data_in(h_col_238), .sum(check_col_238));
bitsadder_128 c_num_239(.data_in(h_col_239), .sum(check_col_239));
bitsadder_128 c_num_240(.data_in(h_col_240), .sum(check_col_240));
bitsadder_128 c_num_241(.data_in(h_col_241), .sum(check_col_241));
bitsadder_128 c_num_242(.data_in(h_col_242), .sum(check_col_242));
bitsadder_128 c_num_243(.data_in(h_col_243), .sum(check_col_243));
bitsadder_128 c_num_244(.data_in(h_col_244), .sum(check_col_244));
bitsadder_128 c_num_245(.data_in(h_col_245), .sum(check_col_245));
bitsadder_128 c_num_246(.data_in(h_col_246), .sum(check_col_246));
bitsadder_128 c_num_247(.data_in(h_col_247), .sum(check_col_247));
bitsadder_128 c_num_248(.data_in(h_col_248), .sum(check_col_248));
bitsadder_128 c_num_249(.data_in(h_col_249), .sum(check_col_249));
bitsadder_128 c_num_250(.data_in(h_col_250), .sum(check_col_250));
bitsadder_128 c_num_251(.data_in(h_col_251), .sum(check_col_251));
bitsadder_128 c_num_252(.data_in(h_col_252), .sum(check_col_252));
bitsadder_128 c_num_253(.data_in(h_col_253), .sum(check_col_253));
bitsadder_128 c_num_254(.data_in(h_col_254), .sum(check_col_254));
bitsadder_128 c_num_255(.data_in(h_col_255), .sum(check_col_255));


bitsadder_128 w_num_0(.data_in(h_col_0 & form_array), .sum(wrong_col_0));
bitsadder_128 w_num_1(.data_in(h_col_1 & form_array), .sum(wrong_col_1));
bitsadder_128 w_num_2(.data_in(h_col_2 & form_array), .sum(wrong_col_2));
bitsadder_128 w_num_3(.data_in(h_col_3 & form_array), .sum(wrong_col_3));
bitsadder_128 w_num_4(.data_in(h_col_4 & form_array), .sum(wrong_col_4));
bitsadder_128 w_num_5(.data_in(h_col_5 & form_array), .sum(wrong_col_5));
bitsadder_128 w_num_6(.data_in(h_col_6 & form_array), .sum(wrong_col_6));
bitsadder_128 w_num_7(.data_in(h_col_7 & form_array), .sum(wrong_col_7));
bitsadder_128 w_num_8(.data_in(h_col_8 & form_array), .sum(wrong_col_8));
bitsadder_128 w_num_9(.data_in(h_col_9 & form_array), .sum(wrong_col_9));
bitsadder_128 w_num_10(.data_in(h_col_10 & form_array), .sum(wrong_col_10));
bitsadder_128 w_num_11(.data_in(h_col_11 & form_array), .sum(wrong_col_11));
bitsadder_128 w_num_12(.data_in(h_col_12 & form_array), .sum(wrong_col_12));
bitsadder_128 w_num_13(.data_in(h_col_13 & form_array), .sum(wrong_col_13));
bitsadder_128 w_num_14(.data_in(h_col_14 & form_array), .sum(wrong_col_14));
bitsadder_128 w_num_15(.data_in(h_col_15 & form_array), .sum(wrong_col_15));
bitsadder_128 w_num_16(.data_in(h_col_16 & form_array), .sum(wrong_col_16));
bitsadder_128 w_num_17(.data_in(h_col_17 & form_array), .sum(wrong_col_17));
bitsadder_128 w_num_18(.data_in(h_col_18 & form_array), .sum(wrong_col_18));
bitsadder_128 w_num_19(.data_in(h_col_19 & form_array), .sum(wrong_col_19));
bitsadder_128 w_num_20(.data_in(h_col_20 & form_array), .sum(wrong_col_20));
bitsadder_128 w_num_21(.data_in(h_col_21 & form_array), .sum(wrong_col_21));
bitsadder_128 w_num_22(.data_in(h_col_22 & form_array), .sum(wrong_col_22));
bitsadder_128 w_num_23(.data_in(h_col_23 & form_array), .sum(wrong_col_23));
bitsadder_128 w_num_24(.data_in(h_col_24 & form_array), .sum(wrong_col_24));
bitsadder_128 w_num_25(.data_in(h_col_25 & form_array), .sum(wrong_col_25));
bitsadder_128 w_num_26(.data_in(h_col_26 & form_array), .sum(wrong_col_26));
bitsadder_128 w_num_27(.data_in(h_col_27 & form_array), .sum(wrong_col_27));
bitsadder_128 w_num_28(.data_in(h_col_28 & form_array), .sum(wrong_col_28));
bitsadder_128 w_num_29(.data_in(h_col_29 & form_array), .sum(wrong_col_29));
bitsadder_128 w_num_30(.data_in(h_col_30 & form_array), .sum(wrong_col_30));
bitsadder_128 w_num_31(.data_in(h_col_31 & form_array), .sum(wrong_col_31));
bitsadder_128 w_num_32(.data_in(h_col_32 & form_array), .sum(wrong_col_32));
bitsadder_128 w_num_33(.data_in(h_col_33 & form_array), .sum(wrong_col_33));
bitsadder_128 w_num_34(.data_in(h_col_34 & form_array), .sum(wrong_col_34));
bitsadder_128 w_num_35(.data_in(h_col_35 & form_array), .sum(wrong_col_35));
bitsadder_128 w_num_36(.data_in(h_col_36 & form_array), .sum(wrong_col_36));
bitsadder_128 w_num_37(.data_in(h_col_37 & form_array), .sum(wrong_col_37));
bitsadder_128 w_num_38(.data_in(h_col_38 & form_array), .sum(wrong_col_38));
bitsadder_128 w_num_39(.data_in(h_col_39 & form_array), .sum(wrong_col_39));
bitsadder_128 w_num_40(.data_in(h_col_40 & form_array), .sum(wrong_col_40));
bitsadder_128 w_num_41(.data_in(h_col_41 & form_array), .sum(wrong_col_41));
bitsadder_128 w_num_42(.data_in(h_col_42 & form_array), .sum(wrong_col_42));
bitsadder_128 w_num_43(.data_in(h_col_43 & form_array), .sum(wrong_col_43));
bitsadder_128 w_num_44(.data_in(h_col_44 & form_array), .sum(wrong_col_44));
bitsadder_128 w_num_45(.data_in(h_col_45 & form_array), .sum(wrong_col_45));
bitsadder_128 w_num_46(.data_in(h_col_46 & form_array), .sum(wrong_col_46));
bitsadder_128 w_num_47(.data_in(h_col_47 & form_array), .sum(wrong_col_47));
bitsadder_128 w_num_48(.data_in(h_col_48 & form_array), .sum(wrong_col_48));
bitsadder_128 w_num_49(.data_in(h_col_49 & form_array), .sum(wrong_col_49));
bitsadder_128 w_num_50(.data_in(h_col_50 & form_array), .sum(wrong_col_50));
bitsadder_128 w_num_51(.data_in(h_col_51 & form_array), .sum(wrong_col_51));
bitsadder_128 w_num_52(.data_in(h_col_52 & form_array), .sum(wrong_col_52));
bitsadder_128 w_num_53(.data_in(h_col_53 & form_array), .sum(wrong_col_53));
bitsadder_128 w_num_54(.data_in(h_col_54 & form_array), .sum(wrong_col_54));
bitsadder_128 w_num_55(.data_in(h_col_55 & form_array), .sum(wrong_col_55));
bitsadder_128 w_num_56(.data_in(h_col_56 & form_array), .sum(wrong_col_56));
bitsadder_128 w_num_57(.data_in(h_col_57 & form_array), .sum(wrong_col_57));
bitsadder_128 w_num_58(.data_in(h_col_58 & form_array), .sum(wrong_col_58));
bitsadder_128 w_num_59(.data_in(h_col_59 & form_array), .sum(wrong_col_59));
bitsadder_128 w_num_60(.data_in(h_col_60 & form_array), .sum(wrong_col_60));
bitsadder_128 w_num_61(.data_in(h_col_61 & form_array), .sum(wrong_col_61));
bitsadder_128 w_num_62(.data_in(h_col_62 & form_array), .sum(wrong_col_62));
bitsadder_128 w_num_63(.data_in(h_col_63 & form_array), .sum(wrong_col_63));
bitsadder_128 w_num_64(.data_in(h_col_64 & form_array), .sum(wrong_col_64));
bitsadder_128 w_num_65(.data_in(h_col_65 & form_array), .sum(wrong_col_65));
bitsadder_128 w_num_66(.data_in(h_col_66 & form_array), .sum(wrong_col_66));
bitsadder_128 w_num_67(.data_in(h_col_67 & form_array), .sum(wrong_col_67));
bitsadder_128 w_num_68(.data_in(h_col_68 & form_array), .sum(wrong_col_68));
bitsadder_128 w_num_69(.data_in(h_col_69 & form_array), .sum(wrong_col_69));
bitsadder_128 w_num_70(.data_in(h_col_70 & form_array), .sum(wrong_col_70));
bitsadder_128 w_num_71(.data_in(h_col_71 & form_array), .sum(wrong_col_71));
bitsadder_128 w_num_72(.data_in(h_col_72 & form_array), .sum(wrong_col_72));
bitsadder_128 w_num_73(.data_in(h_col_73 & form_array), .sum(wrong_col_73));
bitsadder_128 w_num_74(.data_in(h_col_74 & form_array), .sum(wrong_col_74));
bitsadder_128 w_num_75(.data_in(h_col_75 & form_array), .sum(wrong_col_75));
bitsadder_128 w_num_76(.data_in(h_col_76 & form_array), .sum(wrong_col_76));
bitsadder_128 w_num_77(.data_in(h_col_77 & form_array), .sum(wrong_col_77));
bitsadder_128 w_num_78(.data_in(h_col_78 & form_array), .sum(wrong_col_78));
bitsadder_128 w_num_79(.data_in(h_col_79 & form_array), .sum(wrong_col_79));
bitsadder_128 w_num_80(.data_in(h_col_80 & form_array), .sum(wrong_col_80));
bitsadder_128 w_num_81(.data_in(h_col_81 & form_array), .sum(wrong_col_81));
bitsadder_128 w_num_82(.data_in(h_col_82 & form_array), .sum(wrong_col_82));
bitsadder_128 w_num_83(.data_in(h_col_83 & form_array), .sum(wrong_col_83));
bitsadder_128 w_num_84(.data_in(h_col_84 & form_array), .sum(wrong_col_84));
bitsadder_128 w_num_85(.data_in(h_col_85 & form_array), .sum(wrong_col_85));
bitsadder_128 w_num_86(.data_in(h_col_86 & form_array), .sum(wrong_col_86));
bitsadder_128 w_num_87(.data_in(h_col_87 & form_array), .sum(wrong_col_87));
bitsadder_128 w_num_88(.data_in(h_col_88 & form_array), .sum(wrong_col_88));
bitsadder_128 w_num_89(.data_in(h_col_89 & form_array), .sum(wrong_col_89));
bitsadder_128 w_num_90(.data_in(h_col_90 & form_array), .sum(wrong_col_90));
bitsadder_128 w_num_91(.data_in(h_col_91 & form_array), .sum(wrong_col_91));
bitsadder_128 w_num_92(.data_in(h_col_92 & form_array), .sum(wrong_col_92));
bitsadder_128 w_num_93(.data_in(h_col_93 & form_array), .sum(wrong_col_93));
bitsadder_128 w_num_94(.data_in(h_col_94 & form_array), .sum(wrong_col_94));
bitsadder_128 w_num_95(.data_in(h_col_95 & form_array), .sum(wrong_col_95));
bitsadder_128 w_num_96(.data_in(h_col_96 & form_array), .sum(wrong_col_96));
bitsadder_128 w_num_97(.data_in(h_col_97 & form_array), .sum(wrong_col_97));
bitsadder_128 w_num_98(.data_in(h_col_98 & form_array), .sum(wrong_col_98));
bitsadder_128 w_num_99(.data_in(h_col_99 & form_array), .sum(wrong_col_99));
bitsadder_128 w_num_100(.data_in(h_col_100 & form_array), .sum(wrong_col_100));
bitsadder_128 w_num_101(.data_in(h_col_101 & form_array), .sum(wrong_col_101));
bitsadder_128 w_num_102(.data_in(h_col_102 & form_array), .sum(wrong_col_102));
bitsadder_128 w_num_103(.data_in(h_col_103 & form_array), .sum(wrong_col_103));
bitsadder_128 w_num_104(.data_in(h_col_104 & form_array), .sum(wrong_col_104));
bitsadder_128 w_num_105(.data_in(h_col_105 & form_array), .sum(wrong_col_105));
bitsadder_128 w_num_106(.data_in(h_col_106 & form_array), .sum(wrong_col_106));
bitsadder_128 w_num_107(.data_in(h_col_107 & form_array), .sum(wrong_col_107));
bitsadder_128 w_num_108(.data_in(h_col_108 & form_array), .sum(wrong_col_108));
bitsadder_128 w_num_109(.data_in(h_col_109 & form_array), .sum(wrong_col_109));
bitsadder_128 w_num_110(.data_in(h_col_110 & form_array), .sum(wrong_col_110));
bitsadder_128 w_num_111(.data_in(h_col_111 & form_array), .sum(wrong_col_111));
bitsadder_128 w_num_112(.data_in(h_col_112 & form_array), .sum(wrong_col_112));
bitsadder_128 w_num_113(.data_in(h_col_113 & form_array), .sum(wrong_col_113));
bitsadder_128 w_num_114(.data_in(h_col_114 & form_array), .sum(wrong_col_114));
bitsadder_128 w_num_115(.data_in(h_col_115 & form_array), .sum(wrong_col_115));
bitsadder_128 w_num_116(.data_in(h_col_116 & form_array), .sum(wrong_col_116));
bitsadder_128 w_num_117(.data_in(h_col_117 & form_array), .sum(wrong_col_117));
bitsadder_128 w_num_118(.data_in(h_col_118 & form_array), .sum(wrong_col_118));
bitsadder_128 w_num_119(.data_in(h_col_119 & form_array), .sum(wrong_col_119));
bitsadder_128 w_num_120(.data_in(h_col_120 & form_array), .sum(wrong_col_120));
bitsadder_128 w_num_121(.data_in(h_col_121 & form_array), .sum(wrong_col_121));
bitsadder_128 w_num_122(.data_in(h_col_122 & form_array), .sum(wrong_col_122));
bitsadder_128 w_num_123(.data_in(h_col_123 & form_array), .sum(wrong_col_123));
bitsadder_128 w_num_124(.data_in(h_col_124 & form_array), .sum(wrong_col_124));
bitsadder_128 w_num_125(.data_in(h_col_125 & form_array), .sum(wrong_col_125));
bitsadder_128 w_num_126(.data_in(h_col_126 & form_array), .sum(wrong_col_126));
bitsadder_128 w_num_127(.data_in(h_col_127 & form_array), .sum(wrong_col_127));
bitsadder_128 w_num_128(.data_in(h_col_128 & form_array), .sum(wrong_col_128));
bitsadder_128 w_num_129(.data_in(h_col_129 & form_array), .sum(wrong_col_129));
bitsadder_128 w_num_130(.data_in(h_col_130 & form_array), .sum(wrong_col_130));
bitsadder_128 w_num_131(.data_in(h_col_131 & form_array), .sum(wrong_col_131));
bitsadder_128 w_num_132(.data_in(h_col_132 & form_array), .sum(wrong_col_132));
bitsadder_128 w_num_133(.data_in(h_col_133 & form_array), .sum(wrong_col_133));
bitsadder_128 w_num_134(.data_in(h_col_134 & form_array), .sum(wrong_col_134));
bitsadder_128 w_num_135(.data_in(h_col_135 & form_array), .sum(wrong_col_135));
bitsadder_128 w_num_136(.data_in(h_col_136 & form_array), .sum(wrong_col_136));
bitsadder_128 w_num_137(.data_in(h_col_137 & form_array), .sum(wrong_col_137));
bitsadder_128 w_num_138(.data_in(h_col_138 & form_array), .sum(wrong_col_138));
bitsadder_128 w_num_139(.data_in(h_col_139 & form_array), .sum(wrong_col_139));
bitsadder_128 w_num_140(.data_in(h_col_140 & form_array), .sum(wrong_col_140));
bitsadder_128 w_num_141(.data_in(h_col_141 & form_array), .sum(wrong_col_141));
bitsadder_128 w_num_142(.data_in(h_col_142 & form_array), .sum(wrong_col_142));
bitsadder_128 w_num_143(.data_in(h_col_143 & form_array), .sum(wrong_col_143));
bitsadder_128 w_num_144(.data_in(h_col_144 & form_array), .sum(wrong_col_144));
bitsadder_128 w_num_145(.data_in(h_col_145 & form_array), .sum(wrong_col_145));
bitsadder_128 w_num_146(.data_in(h_col_146 & form_array), .sum(wrong_col_146));
bitsadder_128 w_num_147(.data_in(h_col_147 & form_array), .sum(wrong_col_147));
bitsadder_128 w_num_148(.data_in(h_col_148 & form_array), .sum(wrong_col_148));
bitsadder_128 w_num_149(.data_in(h_col_149 & form_array), .sum(wrong_col_149));
bitsadder_128 w_num_150(.data_in(h_col_150 & form_array), .sum(wrong_col_150));
bitsadder_128 w_num_151(.data_in(h_col_151 & form_array), .sum(wrong_col_151));
bitsadder_128 w_num_152(.data_in(h_col_152 & form_array), .sum(wrong_col_152));
bitsadder_128 w_num_153(.data_in(h_col_153 & form_array), .sum(wrong_col_153));
bitsadder_128 w_num_154(.data_in(h_col_154 & form_array), .sum(wrong_col_154));
bitsadder_128 w_num_155(.data_in(h_col_155 & form_array), .sum(wrong_col_155));
bitsadder_128 w_num_156(.data_in(h_col_156 & form_array), .sum(wrong_col_156));
bitsadder_128 w_num_157(.data_in(h_col_157 & form_array), .sum(wrong_col_157));
bitsadder_128 w_num_158(.data_in(h_col_158 & form_array), .sum(wrong_col_158));
bitsadder_128 w_num_159(.data_in(h_col_159 & form_array), .sum(wrong_col_159));
bitsadder_128 w_num_160(.data_in(h_col_160 & form_array), .sum(wrong_col_160));
bitsadder_128 w_num_161(.data_in(h_col_161 & form_array), .sum(wrong_col_161));
bitsadder_128 w_num_162(.data_in(h_col_162 & form_array), .sum(wrong_col_162));
bitsadder_128 w_num_163(.data_in(h_col_163 & form_array), .sum(wrong_col_163));
bitsadder_128 w_num_164(.data_in(h_col_164 & form_array), .sum(wrong_col_164));
bitsadder_128 w_num_165(.data_in(h_col_165 & form_array), .sum(wrong_col_165));
bitsadder_128 w_num_166(.data_in(h_col_166 & form_array), .sum(wrong_col_166));
bitsadder_128 w_num_167(.data_in(h_col_167 & form_array), .sum(wrong_col_167));
bitsadder_128 w_num_168(.data_in(h_col_168 & form_array), .sum(wrong_col_168));
bitsadder_128 w_num_169(.data_in(h_col_169 & form_array), .sum(wrong_col_169));
bitsadder_128 w_num_170(.data_in(h_col_170 & form_array), .sum(wrong_col_170));
bitsadder_128 w_num_171(.data_in(h_col_171 & form_array), .sum(wrong_col_171));
bitsadder_128 w_num_172(.data_in(h_col_172 & form_array), .sum(wrong_col_172));
bitsadder_128 w_num_173(.data_in(h_col_173 & form_array), .sum(wrong_col_173));
bitsadder_128 w_num_174(.data_in(h_col_174 & form_array), .sum(wrong_col_174));
bitsadder_128 w_num_175(.data_in(h_col_175 & form_array), .sum(wrong_col_175));
bitsadder_128 w_num_176(.data_in(h_col_176 & form_array), .sum(wrong_col_176));
bitsadder_128 w_num_177(.data_in(h_col_177 & form_array), .sum(wrong_col_177));
bitsadder_128 w_num_178(.data_in(h_col_178 & form_array), .sum(wrong_col_178));
bitsadder_128 w_num_179(.data_in(h_col_179 & form_array), .sum(wrong_col_179));
bitsadder_128 w_num_180(.data_in(h_col_180 & form_array), .sum(wrong_col_180));
bitsadder_128 w_num_181(.data_in(h_col_181 & form_array), .sum(wrong_col_181));
bitsadder_128 w_num_182(.data_in(h_col_182 & form_array), .sum(wrong_col_182));
bitsadder_128 w_num_183(.data_in(h_col_183 & form_array), .sum(wrong_col_183));
bitsadder_128 w_num_184(.data_in(h_col_184 & form_array), .sum(wrong_col_184));
bitsadder_128 w_num_185(.data_in(h_col_185 & form_array), .sum(wrong_col_185));
bitsadder_128 w_num_186(.data_in(h_col_186 & form_array), .sum(wrong_col_186));
bitsadder_128 w_num_187(.data_in(h_col_187 & form_array), .sum(wrong_col_187));
bitsadder_128 w_num_188(.data_in(h_col_188 & form_array), .sum(wrong_col_188));
bitsadder_128 w_num_189(.data_in(h_col_189 & form_array), .sum(wrong_col_189));
bitsadder_128 w_num_190(.data_in(h_col_190 & form_array), .sum(wrong_col_190));
bitsadder_128 w_num_191(.data_in(h_col_191 & form_array), .sum(wrong_col_191));
bitsadder_128 w_num_192(.data_in(h_col_192 & form_array), .sum(wrong_col_192));
bitsadder_128 w_num_193(.data_in(h_col_193 & form_array), .sum(wrong_col_193));
bitsadder_128 w_num_194(.data_in(h_col_194 & form_array), .sum(wrong_col_194));
bitsadder_128 w_num_195(.data_in(h_col_195 & form_array), .sum(wrong_col_195));
bitsadder_128 w_num_196(.data_in(h_col_196 & form_array), .sum(wrong_col_196));
bitsadder_128 w_num_197(.data_in(h_col_197 & form_array), .sum(wrong_col_197));
bitsadder_128 w_num_198(.data_in(h_col_198 & form_array), .sum(wrong_col_198));
bitsadder_128 w_num_199(.data_in(h_col_199 & form_array), .sum(wrong_col_199));
bitsadder_128 w_num_200(.data_in(h_col_200 & form_array), .sum(wrong_col_200));
bitsadder_128 w_num_201(.data_in(h_col_201 & form_array), .sum(wrong_col_201));
bitsadder_128 w_num_202(.data_in(h_col_202 & form_array), .sum(wrong_col_202));
bitsadder_128 w_num_203(.data_in(h_col_203 & form_array), .sum(wrong_col_203));
bitsadder_128 w_num_204(.data_in(h_col_204 & form_array), .sum(wrong_col_204));
bitsadder_128 w_num_205(.data_in(h_col_205 & form_array), .sum(wrong_col_205));
bitsadder_128 w_num_206(.data_in(h_col_206 & form_array), .sum(wrong_col_206));
bitsadder_128 w_num_207(.data_in(h_col_207 & form_array), .sum(wrong_col_207));
bitsadder_128 w_num_208(.data_in(h_col_208 & form_array), .sum(wrong_col_208));
bitsadder_128 w_num_209(.data_in(h_col_209 & form_array), .sum(wrong_col_209));
bitsadder_128 w_num_210(.data_in(h_col_210 & form_array), .sum(wrong_col_210));
bitsadder_128 w_num_211(.data_in(h_col_211 & form_array), .sum(wrong_col_211));
bitsadder_128 w_num_212(.data_in(h_col_212 & form_array), .sum(wrong_col_212));
bitsadder_128 w_num_213(.data_in(h_col_213 & form_array), .sum(wrong_col_213));
bitsadder_128 w_num_214(.data_in(h_col_214 & form_array), .sum(wrong_col_214));
bitsadder_128 w_num_215(.data_in(h_col_215 & form_array), .sum(wrong_col_215));
bitsadder_128 w_num_216(.data_in(h_col_216 & form_array), .sum(wrong_col_216));
bitsadder_128 w_num_217(.data_in(h_col_217 & form_array), .sum(wrong_col_217));
bitsadder_128 w_num_218(.data_in(h_col_218 & form_array), .sum(wrong_col_218));
bitsadder_128 w_num_219(.data_in(h_col_219 & form_array), .sum(wrong_col_219));
bitsadder_128 w_num_220(.data_in(h_col_220 & form_array), .sum(wrong_col_220));
bitsadder_128 w_num_221(.data_in(h_col_221 & form_array), .sum(wrong_col_221));
bitsadder_128 w_num_222(.data_in(h_col_222 & form_array), .sum(wrong_col_222));
bitsadder_128 w_num_223(.data_in(h_col_223 & form_array), .sum(wrong_col_223));
bitsadder_128 w_num_224(.data_in(h_col_224 & form_array), .sum(wrong_col_224));
bitsadder_128 w_num_225(.data_in(h_col_225 & form_array), .sum(wrong_col_225));
bitsadder_128 w_num_226(.data_in(h_col_226 & form_array), .sum(wrong_col_226));
bitsadder_128 w_num_227(.data_in(h_col_227 & form_array), .sum(wrong_col_227));
bitsadder_128 w_num_228(.data_in(h_col_228 & form_array), .sum(wrong_col_228));
bitsadder_128 w_num_229(.data_in(h_col_229 & form_array), .sum(wrong_col_229));
bitsadder_128 w_num_230(.data_in(h_col_230 & form_array), .sum(wrong_col_230));
bitsadder_128 w_num_231(.data_in(h_col_231 & form_array), .sum(wrong_col_231));
bitsadder_128 w_num_232(.data_in(h_col_232 & form_array), .sum(wrong_col_232));
bitsadder_128 w_num_233(.data_in(h_col_233 & form_array), .sum(wrong_col_233));
bitsadder_128 w_num_234(.data_in(h_col_234 & form_array), .sum(wrong_col_234));
bitsadder_128 w_num_235(.data_in(h_col_235 & form_array), .sum(wrong_col_235));
bitsadder_128 w_num_236(.data_in(h_col_236 & form_array), .sum(wrong_col_236));
bitsadder_128 w_num_237(.data_in(h_col_237 & form_array), .sum(wrong_col_237));
bitsadder_128 w_num_238(.data_in(h_col_238 & form_array), .sum(wrong_col_238));
bitsadder_128 w_num_239(.data_in(h_col_239 & form_array), .sum(wrong_col_239));
bitsadder_128 w_num_240(.data_in(h_col_240 & form_array), .sum(wrong_col_240));
bitsadder_128 w_num_241(.data_in(h_col_241 & form_array), .sum(wrong_col_241));
bitsadder_128 w_num_242(.data_in(h_col_242 & form_array), .sum(wrong_col_242));
bitsadder_128 w_num_243(.data_in(h_col_243 & form_array), .sum(wrong_col_243));
bitsadder_128 w_num_244(.data_in(h_col_244 & form_array), .sum(wrong_col_244));
bitsadder_128 w_num_245(.data_in(h_col_245 & form_array), .sum(wrong_col_245));
bitsadder_128 w_num_246(.data_in(h_col_246 & form_array), .sum(wrong_col_246));
bitsadder_128 w_num_247(.data_in(h_col_247 & form_array), .sum(wrong_col_247));
bitsadder_128 w_num_248(.data_in(h_col_248 & form_array), .sum(wrong_col_248));
bitsadder_128 w_num_249(.data_in(h_col_249 & form_array), .sum(wrong_col_249));
bitsadder_128 w_num_250(.data_in(h_col_250 & form_array), .sum(wrong_col_250));
bitsadder_128 w_num_251(.data_in(h_col_251 & form_array), .sum(wrong_col_251));
bitsadder_128 w_num_252(.data_in(h_col_252 & form_array), .sum(wrong_col_252));
bitsadder_128 w_num_253(.data_in(h_col_253 & form_array), .sum(wrong_col_253));
bitsadder_128 w_num_254(.data_in(h_col_254 & form_array), .sum(wrong_col_254));
bitsadder_128 w_num_255(.data_in(h_col_255 & form_array), .sum(wrong_col_255));


//Edit code:

always@(posedge clk or negedge rst) begin
if(!rst) begin
state <= init;
free_flag <= 1'b0;
valid_flag <= 1'b0;
iter_flag <= 1'b0;
iter_cnt <= 'd0;
deout_reg <= 'd0;
end
else begin

case(state)

init: begin
free_flag <= 1'b1;
tx_buffer <= 'd0;
form_array <= 'd0;
state <= getin;

end


getin: begin
valid_flag <= 1'b0;
if(work) begin
    tx_buffer <= tx;
    update_buffer <= tx;
    form_array <= 'd0;
    free_flag <= 1'b0;
    iter_flag <= 1'b1;
    deout_reg <= 'd0;
    state <= dot;
end
else begin
    if (iter_flag) begin
        tx_buffer <= update_buffer;
        state <= dot;
    end
    else begin
        state <= getin;
    end
end

end


dot: begin

dotarray[0] <= (Harray[0] & tx_buffer);
dotarray[1] <= (Harray[1] & tx_buffer);
dotarray[2] <= (Harray[2] & tx_buffer);
dotarray[3] <= (Harray[3] & tx_buffer);
dotarray[4] <= (Harray[4] & tx_buffer);
dotarray[5] <= (Harray[5] & tx_buffer);
dotarray[6] <= (Harray[6] & tx_buffer);
dotarray[7] <= (Harray[7] & tx_buffer);
dotarray[8] <= (Harray[8] & tx_buffer);
dotarray[9] <= (Harray[9] & tx_buffer);
dotarray[10] <= (Harray[10] & tx_buffer);
dotarray[11] <= (Harray[11] & tx_buffer);
dotarray[12] <= (Harray[12] & tx_buffer);
dotarray[13] <= (Harray[13] & tx_buffer);
dotarray[14] <= (Harray[14] & tx_buffer);
dotarray[15] <= (Harray[15] & tx_buffer);
dotarray[16] <= (Harray[16] & tx_buffer);
dotarray[17] <= (Harray[17] & tx_buffer);
dotarray[18] <= (Harray[18] & tx_buffer);
dotarray[19] <= (Harray[19] & tx_buffer);
dotarray[20] <= (Harray[20] & tx_buffer);
dotarray[21] <= (Harray[21] & tx_buffer);
dotarray[22] <= (Harray[22] & tx_buffer);
dotarray[23] <= (Harray[23] & tx_buffer);
dotarray[24] <= (Harray[24] & tx_buffer);
dotarray[25] <= (Harray[25] & tx_buffer);
dotarray[26] <= (Harray[26] & tx_buffer);
dotarray[27] <= (Harray[27] & tx_buffer);
dotarray[28] <= (Harray[28] & tx_buffer);
dotarray[29] <= (Harray[29] & tx_buffer);
dotarray[30] <= (Harray[30] & tx_buffer);
dotarray[31] <= (Harray[31] & tx_buffer);
dotarray[32] <= (Harray[32] & tx_buffer);
dotarray[33] <= (Harray[33] & tx_buffer);
dotarray[34] <= (Harray[34] & tx_buffer);
dotarray[35] <= (Harray[35] & tx_buffer);
dotarray[36] <= (Harray[36] & tx_buffer);
dotarray[37] <= (Harray[37] & tx_buffer);
dotarray[38] <= (Harray[38] & tx_buffer);
dotarray[39] <= (Harray[39] & tx_buffer);
dotarray[40] <= (Harray[40] & tx_buffer);
dotarray[41] <= (Harray[41] & tx_buffer);
dotarray[42] <= (Harray[42] & tx_buffer);
dotarray[43] <= (Harray[43] & tx_buffer);
dotarray[44] <= (Harray[44] & tx_buffer);
dotarray[45] <= (Harray[45] & tx_buffer);
dotarray[46] <= (Harray[46] & tx_buffer);
dotarray[47] <= (Harray[47] & tx_buffer);
dotarray[48] <= (Harray[48] & tx_buffer);
dotarray[49] <= (Harray[49] & tx_buffer);
dotarray[50] <= (Harray[50] & tx_buffer);
dotarray[51] <= (Harray[51] & tx_buffer);
dotarray[52] <= (Harray[52] & tx_buffer);
dotarray[53] <= (Harray[53] & tx_buffer);
dotarray[54] <= (Harray[54] & tx_buffer);
dotarray[55] <= (Harray[55] & tx_buffer);
dotarray[56] <= (Harray[56] & tx_buffer);
dotarray[57] <= (Harray[57] & tx_buffer);
dotarray[58] <= (Harray[58] & tx_buffer);
dotarray[59] <= (Harray[59] & tx_buffer);
dotarray[60] <= (Harray[60] & tx_buffer);
dotarray[61] <= (Harray[61] & tx_buffer);
dotarray[62] <= (Harray[62] & tx_buffer);
dotarray[63] <= (Harray[63] & tx_buffer);
dotarray[64] <= (Harray[64] & tx_buffer);
dotarray[65] <= (Harray[65] & tx_buffer);
dotarray[66] <= (Harray[66] & tx_buffer);
dotarray[67] <= (Harray[67] & tx_buffer);
dotarray[68] <= (Harray[68] & tx_buffer);
dotarray[69] <= (Harray[69] & tx_buffer);
dotarray[70] <= (Harray[70] & tx_buffer);
dotarray[71] <= (Harray[71] & tx_buffer);
dotarray[72] <= (Harray[72] & tx_buffer);
dotarray[73] <= (Harray[73] & tx_buffer);
dotarray[74] <= (Harray[74] & tx_buffer);
dotarray[75] <= (Harray[75] & tx_buffer);
dotarray[76] <= (Harray[76] & tx_buffer);
dotarray[77] <= (Harray[77] & tx_buffer);
dotarray[78] <= (Harray[78] & tx_buffer);
dotarray[79] <= (Harray[79] & tx_buffer);
dotarray[80] <= (Harray[80] & tx_buffer);
dotarray[81] <= (Harray[81] & tx_buffer);
dotarray[82] <= (Harray[82] & tx_buffer);
dotarray[83] <= (Harray[83] & tx_buffer);
dotarray[84] <= (Harray[84] & tx_buffer);
dotarray[85] <= (Harray[85] & tx_buffer);
dotarray[86] <= (Harray[86] & tx_buffer);
dotarray[87] <= (Harray[87] & tx_buffer);
dotarray[88] <= (Harray[88] & tx_buffer);
dotarray[89] <= (Harray[89] & tx_buffer);
dotarray[90] <= (Harray[90] & tx_buffer);
dotarray[91] <= (Harray[91] & tx_buffer);
dotarray[92] <= (Harray[92] & tx_buffer);
dotarray[93] <= (Harray[93] & tx_buffer);
dotarray[94] <= (Harray[94] & tx_buffer);
dotarray[95] <= (Harray[95] & tx_buffer);
dotarray[96] <= (Harray[96] & tx_buffer);
dotarray[97] <= (Harray[97] & tx_buffer);
dotarray[98] <= (Harray[98] & tx_buffer);
dotarray[99] <= (Harray[99] & tx_buffer);
dotarray[100] <= (Harray[100] & tx_buffer);
dotarray[101] <= (Harray[101] & tx_buffer);
dotarray[102] <= (Harray[102] & tx_buffer);
dotarray[103] <= (Harray[103] & tx_buffer);
dotarray[104] <= (Harray[104] & tx_buffer);
dotarray[105] <= (Harray[105] & tx_buffer);
dotarray[106] <= (Harray[106] & tx_buffer);
dotarray[107] <= (Harray[107] & tx_buffer);
dotarray[108] <= (Harray[108] & tx_buffer);
dotarray[109] <= (Harray[109] & tx_buffer);
dotarray[110] <= (Harray[110] & tx_buffer);
dotarray[111] <= (Harray[111] & tx_buffer);
dotarray[112] <= (Harray[112] & tx_buffer);
dotarray[113] <= (Harray[113] & tx_buffer);
dotarray[114] <= (Harray[114] & tx_buffer);
dotarray[115] <= (Harray[115] & tx_buffer);
dotarray[116] <= (Harray[116] & tx_buffer);
dotarray[117] <= (Harray[117] & tx_buffer);
dotarray[118] <= (Harray[118] & tx_buffer);
dotarray[119] <= (Harray[119] & tx_buffer);
dotarray[120] <= (Harray[120] & tx_buffer);
dotarray[121] <= (Harray[121] & tx_buffer);
dotarray[122] <= (Harray[122] & tx_buffer);
dotarray[123] <= (Harray[123] & tx_buffer);
dotarray[124] <= (Harray[124] & tx_buffer);
dotarray[125] <= (Harray[125] & tx_buffer);
dotarray[126] <= (Harray[126] & tx_buffer);
dotarray[127] <= (Harray[127] & tx_buffer);

state <= judge;

end


judge: begin
form_array <= row_sum_lastbit;
if(row_sum_lastbit == 'd0) begin
    state <= decode;
end
else begin
    valid_flag <= 1'b0;
    state <= check;
end

end


check: begin

check_cnt[0] <= ((check_col_0) >> 1);
check_cnt[1] <= ((check_col_1) >> 1);
check_cnt[2] <= ((check_col_2) >> 1);
check_cnt[3] <= ((check_col_3) >> 1);
check_cnt[4] <= ((check_col_4) >> 1);
check_cnt[5] <= ((check_col_5) >> 1);
check_cnt[6] <= ((check_col_6) >> 1);
check_cnt[7] <= ((check_col_7) >> 1);
check_cnt[8] <= ((check_col_8) >> 1);
check_cnt[9] <= ((check_col_9) >> 1);
check_cnt[10] <= ((check_col_10) >> 1);
check_cnt[11] <= ((check_col_11) >> 1);
check_cnt[12] <= ((check_col_12) >> 1);
check_cnt[13] <= ((check_col_13) >> 1);
check_cnt[14] <= ((check_col_14) >> 1);
check_cnt[15] <= ((check_col_15) >> 1);
check_cnt[16] <= ((check_col_16) >> 1);
check_cnt[17] <= ((check_col_17) >> 1);
check_cnt[18] <= ((check_col_18) >> 1);
check_cnt[19] <= ((check_col_19) >> 1);
check_cnt[20] <= ((check_col_20) >> 1);
check_cnt[21] <= ((check_col_21) >> 1);
check_cnt[22] <= ((check_col_22) >> 1);
check_cnt[23] <= ((check_col_23) >> 1);
check_cnt[24] <= ((check_col_24) >> 1);
check_cnt[25] <= ((check_col_25) >> 1);
check_cnt[26] <= ((check_col_26) >> 1);
check_cnt[27] <= ((check_col_27) >> 1);
check_cnt[28] <= ((check_col_28) >> 1);
check_cnt[29] <= ((check_col_29) >> 1);
check_cnt[30] <= ((check_col_30) >> 1);
check_cnt[31] <= ((check_col_31) >> 1);
check_cnt[32] <= ((check_col_32) >> 1);
check_cnt[33] <= ((check_col_33) >> 1);
check_cnt[34] <= ((check_col_34) >> 1);
check_cnt[35] <= ((check_col_35) >> 1);
check_cnt[36] <= ((check_col_36) >> 1);
check_cnt[37] <= ((check_col_37) >> 1);
check_cnt[38] <= ((check_col_38) >> 1);
check_cnt[39] <= ((check_col_39) >> 1);
check_cnt[40] <= ((check_col_40) >> 1);
check_cnt[41] <= ((check_col_41) >> 1);
check_cnt[42] <= ((check_col_42) >> 1);
check_cnt[43] <= ((check_col_43) >> 1);
check_cnt[44] <= ((check_col_44) >> 1);
check_cnt[45] <= ((check_col_45) >> 1);
check_cnt[46] <= ((check_col_46) >> 1);
check_cnt[47] <= ((check_col_47) >> 1);
check_cnt[48] <= ((check_col_48) >> 1);
check_cnt[49] <= ((check_col_49) >> 1);
check_cnt[50] <= ((check_col_50) >> 1);
check_cnt[51] <= ((check_col_51) >> 1);
check_cnt[52] <= ((check_col_52) >> 1);
check_cnt[53] <= ((check_col_53) >> 1);
check_cnt[54] <= ((check_col_54) >> 1);
check_cnt[55] <= ((check_col_55) >> 1);
check_cnt[56] <= ((check_col_56) >> 1);
check_cnt[57] <= ((check_col_57) >> 1);
check_cnt[58] <= ((check_col_58) >> 1);
check_cnt[59] <= ((check_col_59) >> 1);
check_cnt[60] <= ((check_col_60) >> 1);
check_cnt[61] <= ((check_col_61) >> 1);
check_cnt[62] <= ((check_col_62) >> 1);
check_cnt[63] <= ((check_col_63) >> 1);
check_cnt[64] <= ((check_col_64) >> 1);
check_cnt[65] <= ((check_col_65) >> 1);
check_cnt[66] <= ((check_col_66) >> 1);
check_cnt[67] <= ((check_col_67) >> 1);
check_cnt[68] <= ((check_col_68) >> 1);
check_cnt[69] <= ((check_col_69) >> 1);
check_cnt[70] <= ((check_col_70) >> 1);
check_cnt[71] <= ((check_col_71) >> 1);
check_cnt[72] <= ((check_col_72) >> 1);
check_cnt[73] <= ((check_col_73) >> 1);
check_cnt[74] <= ((check_col_74) >> 1);
check_cnt[75] <= ((check_col_75) >> 1);
check_cnt[76] <= ((check_col_76) >> 1);
check_cnt[77] <= ((check_col_77) >> 1);
check_cnt[78] <= ((check_col_78) >> 1);
check_cnt[79] <= ((check_col_79) >> 1);
check_cnt[80] <= ((check_col_80) >> 1);
check_cnt[81] <= ((check_col_81) >> 1);
check_cnt[82] <= ((check_col_82) >> 1);
check_cnt[83] <= ((check_col_83) >> 1);
check_cnt[84] <= ((check_col_84) >> 1);
check_cnt[85] <= ((check_col_85) >> 1);
check_cnt[86] <= ((check_col_86) >> 1);
check_cnt[87] <= ((check_col_87) >> 1);
check_cnt[88] <= ((check_col_88) >> 1);
check_cnt[89] <= ((check_col_89) >> 1);
check_cnt[90] <= ((check_col_90) >> 1);
check_cnt[91] <= ((check_col_91) >> 1);
check_cnt[92] <= ((check_col_92) >> 1);
check_cnt[93] <= ((check_col_93) >> 1);
check_cnt[94] <= ((check_col_94) >> 1);
check_cnt[95] <= ((check_col_95) >> 1);
check_cnt[96] <= ((check_col_96) >> 1);
check_cnt[97] <= ((check_col_97) >> 1);
check_cnt[98] <= ((check_col_98) >> 1);
check_cnt[99] <= ((check_col_99) >> 1);
check_cnt[100] <= ((check_col_100) >> 1);
check_cnt[101] <= ((check_col_101) >> 1);
check_cnt[102] <= ((check_col_102) >> 1);
check_cnt[103] <= ((check_col_103) >> 1);
check_cnt[104] <= ((check_col_104) >> 1);
check_cnt[105] <= ((check_col_105) >> 1);
check_cnt[106] <= ((check_col_106) >> 1);
check_cnt[107] <= ((check_col_107) >> 1);
check_cnt[108] <= ((check_col_108) >> 1);
check_cnt[109] <= ((check_col_109) >> 1);
check_cnt[110] <= ((check_col_110) >> 1);
check_cnt[111] <= ((check_col_111) >> 1);
check_cnt[112] <= ((check_col_112) >> 1);
check_cnt[113] <= ((check_col_113) >> 1);
check_cnt[114] <= ((check_col_114) >> 1);
check_cnt[115] <= ((check_col_115) >> 1);
check_cnt[116] <= ((check_col_116) >> 1);
check_cnt[117] <= ((check_col_117) >> 1);
check_cnt[118] <= ((check_col_118) >> 1);
check_cnt[119] <= ((check_col_119) >> 1);
check_cnt[120] <= ((check_col_120) >> 1);
check_cnt[121] <= ((check_col_121) >> 1);
check_cnt[122] <= ((check_col_122) >> 1);
check_cnt[123] <= ((check_col_123) >> 1);
check_cnt[124] <= ((check_col_124) >> 1);
check_cnt[125] <= ((check_col_125) >> 1);
check_cnt[126] <= ((check_col_126) >> 1);
check_cnt[127] <= ((check_col_127) >> 1);
check_cnt[128] <= ((check_col_128) >> 1);
check_cnt[129] <= ((check_col_129) >> 1);
check_cnt[130] <= ((check_col_130) >> 1);
check_cnt[131] <= ((check_col_131) >> 1);
check_cnt[132] <= ((check_col_132) >> 1);
check_cnt[133] <= ((check_col_133) >> 1);
check_cnt[134] <= ((check_col_134) >> 1);
check_cnt[135] <= ((check_col_135) >> 1);
check_cnt[136] <= ((check_col_136) >> 1);
check_cnt[137] <= ((check_col_137) >> 1);
check_cnt[138] <= ((check_col_138) >> 1);
check_cnt[139] <= ((check_col_139) >> 1);
check_cnt[140] <= ((check_col_140) >> 1);
check_cnt[141] <= ((check_col_141) >> 1);
check_cnt[142] <= ((check_col_142) >> 1);
check_cnt[143] <= ((check_col_143) >> 1);
check_cnt[144] <= ((check_col_144) >> 1);
check_cnt[145] <= ((check_col_145) >> 1);
check_cnt[146] <= ((check_col_146) >> 1);
check_cnt[147] <= ((check_col_147) >> 1);
check_cnt[148] <= ((check_col_148) >> 1);
check_cnt[149] <= ((check_col_149) >> 1);
check_cnt[150] <= ((check_col_150) >> 1);
check_cnt[151] <= ((check_col_151) >> 1);
check_cnt[152] <= ((check_col_152) >> 1);
check_cnt[153] <= ((check_col_153) >> 1);
check_cnt[154] <= ((check_col_154) >> 1);
check_cnt[155] <= ((check_col_155) >> 1);
check_cnt[156] <= ((check_col_156) >> 1);
check_cnt[157] <= ((check_col_157) >> 1);
check_cnt[158] <= ((check_col_158) >> 1);
check_cnt[159] <= ((check_col_159) >> 1);
check_cnt[160] <= ((check_col_160) >> 1);
check_cnt[161] <= ((check_col_161) >> 1);
check_cnt[162] <= ((check_col_162) >> 1);
check_cnt[163] <= ((check_col_163) >> 1);
check_cnt[164] <= ((check_col_164) >> 1);
check_cnt[165] <= ((check_col_165) >> 1);
check_cnt[166] <= ((check_col_166) >> 1);
check_cnt[167] <= ((check_col_167) >> 1);
check_cnt[168] <= ((check_col_168) >> 1);
check_cnt[169] <= ((check_col_169) >> 1);
check_cnt[170] <= ((check_col_170) >> 1);
check_cnt[171] <= ((check_col_171) >> 1);
check_cnt[172] <= ((check_col_172) >> 1);
check_cnt[173] <= ((check_col_173) >> 1);
check_cnt[174] <= ((check_col_174) >> 1);
check_cnt[175] <= ((check_col_175) >> 1);
check_cnt[176] <= ((check_col_176) >> 1);
check_cnt[177] <= ((check_col_177) >> 1);
check_cnt[178] <= ((check_col_178) >> 1);
check_cnt[179] <= ((check_col_179) >> 1);
check_cnt[180] <= ((check_col_180) >> 1);
check_cnt[181] <= ((check_col_181) >> 1);
check_cnt[182] <= ((check_col_182) >> 1);
check_cnt[183] <= ((check_col_183) >> 1);
check_cnt[184] <= ((check_col_184) >> 1);
check_cnt[185] <= ((check_col_185) >> 1);
check_cnt[186] <= ((check_col_186) >> 1);
check_cnt[187] <= ((check_col_187) >> 1);
check_cnt[188] <= ((check_col_188) >> 1);
check_cnt[189] <= ((check_col_189) >> 1);
check_cnt[190] <= ((check_col_190) >> 1);
check_cnt[191] <= ((check_col_191) >> 1);
check_cnt[192] <= ((check_col_192) >> 1);
check_cnt[193] <= ((check_col_193) >> 1);
check_cnt[194] <= ((check_col_194) >> 1);
check_cnt[195] <= ((check_col_195) >> 1);
check_cnt[196] <= ((check_col_196) >> 1);
check_cnt[197] <= ((check_col_197) >> 1);
check_cnt[198] <= ((check_col_198) >> 1);
check_cnt[199] <= ((check_col_199) >> 1);
check_cnt[200] <= ((check_col_200) >> 1);
check_cnt[201] <= ((check_col_201) >> 1);
check_cnt[202] <= ((check_col_202) >> 1);
check_cnt[203] <= ((check_col_203) >> 1);
check_cnt[204] <= ((check_col_204) >> 1);
check_cnt[205] <= ((check_col_205) >> 1);
check_cnt[206] <= ((check_col_206) >> 1);
check_cnt[207] <= ((check_col_207) >> 1);
check_cnt[208] <= ((check_col_208) >> 1);
check_cnt[209] <= ((check_col_209) >> 1);
check_cnt[210] <= ((check_col_210) >> 1);
check_cnt[211] <= ((check_col_211) >> 1);
check_cnt[212] <= ((check_col_212) >> 1);
check_cnt[213] <= ((check_col_213) >> 1);
check_cnt[214] <= ((check_col_214) >> 1);
check_cnt[215] <= ((check_col_215) >> 1);
check_cnt[216] <= ((check_col_216) >> 1);
check_cnt[217] <= ((check_col_217) >> 1);
check_cnt[218] <= ((check_col_218) >> 1);
check_cnt[219] <= ((check_col_219) >> 1);
check_cnt[220] <= ((check_col_220) >> 1);
check_cnt[221] <= ((check_col_221) >> 1);
check_cnt[222] <= ((check_col_222) >> 1);
check_cnt[223] <= ((check_col_223) >> 1);
check_cnt[224] <= ((check_col_224) >> 1);
check_cnt[225] <= ((check_col_225) >> 1);
check_cnt[226] <= ((check_col_226) >> 1);
check_cnt[227] <= ((check_col_227) >> 1);
check_cnt[228] <= ((check_col_228) >> 1);
check_cnt[229] <= ((check_col_229) >> 1);
check_cnt[230] <= ((check_col_230) >> 1);
check_cnt[231] <= ((check_col_231) >> 1);
check_cnt[232] <= ((check_col_232) >> 1);
check_cnt[233] <= ((check_col_233) >> 1);
check_cnt[234] <= ((check_col_234) >> 1);
check_cnt[235] <= ((check_col_235) >> 1);
check_cnt[236] <= ((check_col_236) >> 1);
check_cnt[237] <= ((check_col_237) >> 1);
check_cnt[238] <= ((check_col_238) >> 1);
check_cnt[239] <= ((check_col_239) >> 1);
check_cnt[240] <= ((check_col_240) >> 1);
check_cnt[241] <= ((check_col_241) >> 1);
check_cnt[242] <= ((check_col_242) >> 1);
check_cnt[243] <= ((check_col_243) >> 1);
check_cnt[244] <= ((check_col_244) >> 1);
check_cnt[245] <= ((check_col_245) >> 1);
check_cnt[246] <= ((check_col_246) >> 1);
check_cnt[247] <= ((check_col_247) >> 1);
check_cnt[248] <= ((check_col_248) >> 1);
check_cnt[249] <= ((check_col_249) >> 1);
check_cnt[250] <= ((check_col_250) >> 1);
check_cnt[251] <= ((check_col_251) >> 1);
check_cnt[252] <= ((check_col_252) >> 1);
check_cnt[253] <= ((check_col_253) >> 1);
check_cnt[254] <= ((check_col_254) >> 1);
check_cnt[255] <= ((check_col_255) >> 1);

wrong_cnt[0] <= wrong_col_0;
wrong_cnt[1] <= wrong_col_1;
wrong_cnt[2] <= wrong_col_2;
wrong_cnt[3] <= wrong_col_3;
wrong_cnt[4] <= wrong_col_4;
wrong_cnt[5] <= wrong_col_5;
wrong_cnt[6] <= wrong_col_6;
wrong_cnt[7] <= wrong_col_7;
wrong_cnt[8] <= wrong_col_8;
wrong_cnt[9] <= wrong_col_9;
wrong_cnt[10] <= wrong_col_10;
wrong_cnt[11] <= wrong_col_11;
wrong_cnt[12] <= wrong_col_12;
wrong_cnt[13] <= wrong_col_13;
wrong_cnt[14] <= wrong_col_14;
wrong_cnt[15] <= wrong_col_15;
wrong_cnt[16] <= wrong_col_16;
wrong_cnt[17] <= wrong_col_17;
wrong_cnt[18] <= wrong_col_18;
wrong_cnt[19] <= wrong_col_19;
wrong_cnt[20] <= wrong_col_20;
wrong_cnt[21] <= wrong_col_21;
wrong_cnt[22] <= wrong_col_22;
wrong_cnt[23] <= wrong_col_23;
wrong_cnt[24] <= wrong_col_24;
wrong_cnt[25] <= wrong_col_25;
wrong_cnt[26] <= wrong_col_26;
wrong_cnt[27] <= wrong_col_27;
wrong_cnt[28] <= wrong_col_28;
wrong_cnt[29] <= wrong_col_29;
wrong_cnt[30] <= wrong_col_30;
wrong_cnt[31] <= wrong_col_31;
wrong_cnt[32] <= wrong_col_32;
wrong_cnt[33] <= wrong_col_33;
wrong_cnt[34] <= wrong_col_34;
wrong_cnt[35] <= wrong_col_35;
wrong_cnt[36] <= wrong_col_36;
wrong_cnt[37] <= wrong_col_37;
wrong_cnt[38] <= wrong_col_38;
wrong_cnt[39] <= wrong_col_39;
wrong_cnt[40] <= wrong_col_40;
wrong_cnt[41] <= wrong_col_41;
wrong_cnt[42] <= wrong_col_42;
wrong_cnt[43] <= wrong_col_43;
wrong_cnt[44] <= wrong_col_44;
wrong_cnt[45] <= wrong_col_45;
wrong_cnt[46] <= wrong_col_46;
wrong_cnt[47] <= wrong_col_47;
wrong_cnt[48] <= wrong_col_48;
wrong_cnt[49] <= wrong_col_49;
wrong_cnt[50] <= wrong_col_50;
wrong_cnt[51] <= wrong_col_51;
wrong_cnt[52] <= wrong_col_52;
wrong_cnt[53] <= wrong_col_53;
wrong_cnt[54] <= wrong_col_54;
wrong_cnt[55] <= wrong_col_55;
wrong_cnt[56] <= wrong_col_56;
wrong_cnt[57] <= wrong_col_57;
wrong_cnt[58] <= wrong_col_58;
wrong_cnt[59] <= wrong_col_59;
wrong_cnt[60] <= wrong_col_60;
wrong_cnt[61] <= wrong_col_61;
wrong_cnt[62] <= wrong_col_62;
wrong_cnt[63] <= wrong_col_63;
wrong_cnt[64] <= wrong_col_64;
wrong_cnt[65] <= wrong_col_65;
wrong_cnt[66] <= wrong_col_66;
wrong_cnt[67] <= wrong_col_67;
wrong_cnt[68] <= wrong_col_68;
wrong_cnt[69] <= wrong_col_69;
wrong_cnt[70] <= wrong_col_70;
wrong_cnt[71] <= wrong_col_71;
wrong_cnt[72] <= wrong_col_72;
wrong_cnt[73] <= wrong_col_73;
wrong_cnt[74] <= wrong_col_74;
wrong_cnt[75] <= wrong_col_75;
wrong_cnt[76] <= wrong_col_76;
wrong_cnt[77] <= wrong_col_77;
wrong_cnt[78] <= wrong_col_78;
wrong_cnt[79] <= wrong_col_79;
wrong_cnt[80] <= wrong_col_80;
wrong_cnt[81] <= wrong_col_81;
wrong_cnt[82] <= wrong_col_82;
wrong_cnt[83] <= wrong_col_83;
wrong_cnt[84] <= wrong_col_84;
wrong_cnt[85] <= wrong_col_85;
wrong_cnt[86] <= wrong_col_86;
wrong_cnt[87] <= wrong_col_87;
wrong_cnt[88] <= wrong_col_88;
wrong_cnt[89] <= wrong_col_89;
wrong_cnt[90] <= wrong_col_90;
wrong_cnt[91] <= wrong_col_91;
wrong_cnt[92] <= wrong_col_92;
wrong_cnt[93] <= wrong_col_93;
wrong_cnt[94] <= wrong_col_94;
wrong_cnt[95] <= wrong_col_95;
wrong_cnt[96] <= wrong_col_96;
wrong_cnt[97] <= wrong_col_97;
wrong_cnt[98] <= wrong_col_98;
wrong_cnt[99] <= wrong_col_99;
wrong_cnt[100] <= wrong_col_100;
wrong_cnt[101] <= wrong_col_101;
wrong_cnt[102] <= wrong_col_102;
wrong_cnt[103] <= wrong_col_103;
wrong_cnt[104] <= wrong_col_104;
wrong_cnt[105] <= wrong_col_105;
wrong_cnt[106] <= wrong_col_106;
wrong_cnt[107] <= wrong_col_107;
wrong_cnt[108] <= wrong_col_108;
wrong_cnt[109] <= wrong_col_109;
wrong_cnt[110] <= wrong_col_110;
wrong_cnt[111] <= wrong_col_111;
wrong_cnt[112] <= wrong_col_112;
wrong_cnt[113] <= wrong_col_113;
wrong_cnt[114] <= wrong_col_114;
wrong_cnt[115] <= wrong_col_115;
wrong_cnt[116] <= wrong_col_116;
wrong_cnt[117] <= wrong_col_117;
wrong_cnt[118] <= wrong_col_118;
wrong_cnt[119] <= wrong_col_119;
wrong_cnt[120] <= wrong_col_120;
wrong_cnt[121] <= wrong_col_121;
wrong_cnt[122] <= wrong_col_122;
wrong_cnt[123] <= wrong_col_123;
wrong_cnt[124] <= wrong_col_124;
wrong_cnt[125] <= wrong_col_125;
wrong_cnt[126] <= wrong_col_126;
wrong_cnt[127] <= wrong_col_127;
wrong_cnt[128] <= wrong_col_128;
wrong_cnt[129] <= wrong_col_129;
wrong_cnt[130] <= wrong_col_130;
wrong_cnt[131] <= wrong_col_131;
wrong_cnt[132] <= wrong_col_132;
wrong_cnt[133] <= wrong_col_133;
wrong_cnt[134] <= wrong_col_134;
wrong_cnt[135] <= wrong_col_135;
wrong_cnt[136] <= wrong_col_136;
wrong_cnt[137] <= wrong_col_137;
wrong_cnt[138] <= wrong_col_138;
wrong_cnt[139] <= wrong_col_139;
wrong_cnt[140] <= wrong_col_140;
wrong_cnt[141] <= wrong_col_141;
wrong_cnt[142] <= wrong_col_142;
wrong_cnt[143] <= wrong_col_143;
wrong_cnt[144] <= wrong_col_144;
wrong_cnt[145] <= wrong_col_145;
wrong_cnt[146] <= wrong_col_146;
wrong_cnt[147] <= wrong_col_147;
wrong_cnt[148] <= wrong_col_148;
wrong_cnt[149] <= wrong_col_149;
wrong_cnt[150] <= wrong_col_150;
wrong_cnt[151] <= wrong_col_151;
wrong_cnt[152] <= wrong_col_152;
wrong_cnt[153] <= wrong_col_153;
wrong_cnt[154] <= wrong_col_154;
wrong_cnt[155] <= wrong_col_155;
wrong_cnt[156] <= wrong_col_156;
wrong_cnt[157] <= wrong_col_157;
wrong_cnt[158] <= wrong_col_158;
wrong_cnt[159] <= wrong_col_159;
wrong_cnt[160] <= wrong_col_160;
wrong_cnt[161] <= wrong_col_161;
wrong_cnt[162] <= wrong_col_162;
wrong_cnt[163] <= wrong_col_163;
wrong_cnt[164] <= wrong_col_164;
wrong_cnt[165] <= wrong_col_165;
wrong_cnt[166] <= wrong_col_166;
wrong_cnt[167] <= wrong_col_167;
wrong_cnt[168] <= wrong_col_168;
wrong_cnt[169] <= wrong_col_169;
wrong_cnt[170] <= wrong_col_170;
wrong_cnt[171] <= wrong_col_171;
wrong_cnt[172] <= wrong_col_172;
wrong_cnt[173] <= wrong_col_173;
wrong_cnt[174] <= wrong_col_174;
wrong_cnt[175] <= wrong_col_175;
wrong_cnt[176] <= wrong_col_176;
wrong_cnt[177] <= wrong_col_177;
wrong_cnt[178] <= wrong_col_178;
wrong_cnt[179] <= wrong_col_179;
wrong_cnt[180] <= wrong_col_180;
wrong_cnt[181] <= wrong_col_181;
wrong_cnt[182] <= wrong_col_182;
wrong_cnt[183] <= wrong_col_183;
wrong_cnt[184] <= wrong_col_184;
wrong_cnt[185] <= wrong_col_185;
wrong_cnt[186] <= wrong_col_186;
wrong_cnt[187] <= wrong_col_187;
wrong_cnt[188] <= wrong_col_188;
wrong_cnt[189] <= wrong_col_189;
wrong_cnt[190] <= wrong_col_190;
wrong_cnt[191] <= wrong_col_191;
wrong_cnt[192] <= wrong_col_192;
wrong_cnt[193] <= wrong_col_193;
wrong_cnt[194] <= wrong_col_194;
wrong_cnt[195] <= wrong_col_195;
wrong_cnt[196] <= wrong_col_196;
wrong_cnt[197] <= wrong_col_197;
wrong_cnt[198] <= wrong_col_198;
wrong_cnt[199] <= wrong_col_199;
wrong_cnt[200] <= wrong_col_200;
wrong_cnt[201] <= wrong_col_201;
wrong_cnt[202] <= wrong_col_202;
wrong_cnt[203] <= wrong_col_203;
wrong_cnt[204] <= wrong_col_204;
wrong_cnt[205] <= wrong_col_205;
wrong_cnt[206] <= wrong_col_206;
wrong_cnt[207] <= wrong_col_207;
wrong_cnt[208] <= wrong_col_208;
wrong_cnt[209] <= wrong_col_209;
wrong_cnt[210] <= wrong_col_210;
wrong_cnt[211] <= wrong_col_211;
wrong_cnt[212] <= wrong_col_212;
wrong_cnt[213] <= wrong_col_213;
wrong_cnt[214] <= wrong_col_214;
wrong_cnt[215] <= wrong_col_215;
wrong_cnt[216] <= wrong_col_216;
wrong_cnt[217] <= wrong_col_217;
wrong_cnt[218] <= wrong_col_218;
wrong_cnt[219] <= wrong_col_219;
wrong_cnt[220] <= wrong_col_220;
wrong_cnt[221] <= wrong_col_221;
wrong_cnt[222] <= wrong_col_222;
wrong_cnt[223] <= wrong_col_223;
wrong_cnt[224] <= wrong_col_224;
wrong_cnt[225] <= wrong_col_225;
wrong_cnt[226] <= wrong_col_226;
wrong_cnt[227] <= wrong_col_227;
wrong_cnt[228] <= wrong_col_228;
wrong_cnt[229] <= wrong_col_229;
wrong_cnt[230] <= wrong_col_230;
wrong_cnt[231] <= wrong_col_231;
wrong_cnt[232] <= wrong_col_232;
wrong_cnt[233] <= wrong_col_233;
wrong_cnt[234] <= wrong_col_234;
wrong_cnt[235] <= wrong_col_235;
wrong_cnt[236] <= wrong_col_236;
wrong_cnt[237] <= wrong_col_237;
wrong_cnt[238] <= wrong_col_238;
wrong_cnt[239] <= wrong_col_239;
wrong_cnt[240] <= wrong_col_240;
wrong_cnt[241] <= wrong_col_241;
wrong_cnt[242] <= wrong_col_242;
wrong_cnt[243] <= wrong_col_243;
wrong_cnt[244] <= wrong_col_244;
wrong_cnt[245] <= wrong_col_245;
wrong_cnt[246] <= wrong_col_246;
wrong_cnt[247] <= wrong_col_247;
wrong_cnt[248] <= wrong_col_248;
wrong_cnt[249] <= wrong_col_249;
wrong_cnt[250] <= wrong_col_250;
wrong_cnt[251] <= wrong_col_251;
wrong_cnt[252] <= wrong_col_252;
wrong_cnt[253] <= wrong_col_253;
wrong_cnt[254] <= wrong_col_254;
wrong_cnt[255] <= wrong_col_255;

state <= compare;

end


compare: begin

if(wrong_cnt[0] > check_cnt[0]) begin update_buffer[0] <= ~tx_buffer[0]; end else begin update_buffer[0] <= tx_buffer[0]; end
if(wrong_cnt[1] > check_cnt[1]) begin update_buffer[1] <= ~tx_buffer[1]; end else begin update_buffer[1] <= tx_buffer[1]; end
if(wrong_cnt[2] > check_cnt[2]) begin update_buffer[2] <= ~tx_buffer[2]; end else begin update_buffer[2] <= tx_buffer[2]; end
if(wrong_cnt[3] > check_cnt[3]) begin update_buffer[3] <= ~tx_buffer[3]; end else begin update_buffer[3] <= tx_buffer[3]; end
if(wrong_cnt[4] > check_cnt[4]) begin update_buffer[4] <= ~tx_buffer[4]; end else begin update_buffer[4] <= tx_buffer[4]; end
if(wrong_cnt[5] > check_cnt[5]) begin update_buffer[5] <= ~tx_buffer[5]; end else begin update_buffer[5] <= tx_buffer[5]; end
if(wrong_cnt[6] > check_cnt[6]) begin update_buffer[6] <= ~tx_buffer[6]; end else begin update_buffer[6] <= tx_buffer[6]; end
if(wrong_cnt[7] > check_cnt[7]) begin update_buffer[7] <= ~tx_buffer[7]; end else begin update_buffer[7] <= tx_buffer[7]; end
if(wrong_cnt[8] > check_cnt[8]) begin update_buffer[8] <= ~tx_buffer[8]; end else begin update_buffer[8] <= tx_buffer[8]; end
if(wrong_cnt[9] > check_cnt[9]) begin update_buffer[9] <= ~tx_buffer[9]; end else begin update_buffer[9] <= tx_buffer[9]; end
if(wrong_cnt[10] > check_cnt[10]) begin update_buffer[10] <= ~tx_buffer[10]; end else begin update_buffer[10] <= tx_buffer[10]; end
if(wrong_cnt[11] > check_cnt[11]) begin update_buffer[11] <= ~tx_buffer[11]; end else begin update_buffer[11] <= tx_buffer[11]; end
if(wrong_cnt[12] > check_cnt[12]) begin update_buffer[12] <= ~tx_buffer[12]; end else begin update_buffer[12] <= tx_buffer[12]; end
if(wrong_cnt[13] > check_cnt[13]) begin update_buffer[13] <= ~tx_buffer[13]; end else begin update_buffer[13] <= tx_buffer[13]; end
if(wrong_cnt[14] > check_cnt[14]) begin update_buffer[14] <= ~tx_buffer[14]; end else begin update_buffer[14] <= tx_buffer[14]; end
if(wrong_cnt[15] > check_cnt[15]) begin update_buffer[15] <= ~tx_buffer[15]; end else begin update_buffer[15] <= tx_buffer[15]; end
if(wrong_cnt[16] > check_cnt[16]) begin update_buffer[16] <= ~tx_buffer[16]; end else begin update_buffer[16] <= tx_buffer[16]; end
if(wrong_cnt[17] > check_cnt[17]) begin update_buffer[17] <= ~tx_buffer[17]; end else begin update_buffer[17] <= tx_buffer[17]; end
if(wrong_cnt[18] > check_cnt[18]) begin update_buffer[18] <= ~tx_buffer[18]; end else begin update_buffer[18] <= tx_buffer[18]; end
if(wrong_cnt[19] > check_cnt[19]) begin update_buffer[19] <= ~tx_buffer[19]; end else begin update_buffer[19] <= tx_buffer[19]; end
if(wrong_cnt[20] > check_cnt[20]) begin update_buffer[20] <= ~tx_buffer[20]; end else begin update_buffer[20] <= tx_buffer[20]; end
if(wrong_cnt[21] > check_cnt[21]) begin update_buffer[21] <= ~tx_buffer[21]; end else begin update_buffer[21] <= tx_buffer[21]; end
if(wrong_cnt[22] > check_cnt[22]) begin update_buffer[22] <= ~tx_buffer[22]; end else begin update_buffer[22] <= tx_buffer[22]; end
if(wrong_cnt[23] > check_cnt[23]) begin update_buffer[23] <= ~tx_buffer[23]; end else begin update_buffer[23] <= tx_buffer[23]; end
if(wrong_cnt[24] > check_cnt[24]) begin update_buffer[24] <= ~tx_buffer[24]; end else begin update_buffer[24] <= tx_buffer[24]; end
if(wrong_cnt[25] > check_cnt[25]) begin update_buffer[25] <= ~tx_buffer[25]; end else begin update_buffer[25] <= tx_buffer[25]; end
if(wrong_cnt[26] > check_cnt[26]) begin update_buffer[26] <= ~tx_buffer[26]; end else begin update_buffer[26] <= tx_buffer[26]; end
if(wrong_cnt[27] > check_cnt[27]) begin update_buffer[27] <= ~tx_buffer[27]; end else begin update_buffer[27] <= tx_buffer[27]; end
if(wrong_cnt[28] > check_cnt[28]) begin update_buffer[28] <= ~tx_buffer[28]; end else begin update_buffer[28] <= tx_buffer[28]; end
if(wrong_cnt[29] > check_cnt[29]) begin update_buffer[29] <= ~tx_buffer[29]; end else begin update_buffer[29] <= tx_buffer[29]; end
if(wrong_cnt[30] > check_cnt[30]) begin update_buffer[30] <= ~tx_buffer[30]; end else begin update_buffer[30] <= tx_buffer[30]; end
if(wrong_cnt[31] > check_cnt[31]) begin update_buffer[31] <= ~tx_buffer[31]; end else begin update_buffer[31] <= tx_buffer[31]; end
if(wrong_cnt[32] > check_cnt[32]) begin update_buffer[32] <= ~tx_buffer[32]; end else begin update_buffer[32] <= tx_buffer[32]; end
if(wrong_cnt[33] > check_cnt[33]) begin update_buffer[33] <= ~tx_buffer[33]; end else begin update_buffer[33] <= tx_buffer[33]; end
if(wrong_cnt[34] > check_cnt[34]) begin update_buffer[34] <= ~tx_buffer[34]; end else begin update_buffer[34] <= tx_buffer[34]; end
if(wrong_cnt[35] > check_cnt[35]) begin update_buffer[35] <= ~tx_buffer[35]; end else begin update_buffer[35] <= tx_buffer[35]; end
if(wrong_cnt[36] > check_cnt[36]) begin update_buffer[36] <= ~tx_buffer[36]; end else begin update_buffer[36] <= tx_buffer[36]; end
if(wrong_cnt[37] > check_cnt[37]) begin update_buffer[37] <= ~tx_buffer[37]; end else begin update_buffer[37] <= tx_buffer[37]; end
if(wrong_cnt[38] > check_cnt[38]) begin update_buffer[38] <= ~tx_buffer[38]; end else begin update_buffer[38] <= tx_buffer[38]; end
if(wrong_cnt[39] > check_cnt[39]) begin update_buffer[39] <= ~tx_buffer[39]; end else begin update_buffer[39] <= tx_buffer[39]; end
if(wrong_cnt[40] > check_cnt[40]) begin update_buffer[40] <= ~tx_buffer[40]; end else begin update_buffer[40] <= tx_buffer[40]; end
if(wrong_cnt[41] > check_cnt[41]) begin update_buffer[41] <= ~tx_buffer[41]; end else begin update_buffer[41] <= tx_buffer[41]; end
if(wrong_cnt[42] > check_cnt[42]) begin update_buffer[42] <= ~tx_buffer[42]; end else begin update_buffer[42] <= tx_buffer[42]; end
if(wrong_cnt[43] > check_cnt[43]) begin update_buffer[43] <= ~tx_buffer[43]; end else begin update_buffer[43] <= tx_buffer[43]; end
if(wrong_cnt[44] > check_cnt[44]) begin update_buffer[44] <= ~tx_buffer[44]; end else begin update_buffer[44] <= tx_buffer[44]; end
if(wrong_cnt[45] > check_cnt[45]) begin update_buffer[45] <= ~tx_buffer[45]; end else begin update_buffer[45] <= tx_buffer[45]; end
if(wrong_cnt[46] > check_cnt[46]) begin update_buffer[46] <= ~tx_buffer[46]; end else begin update_buffer[46] <= tx_buffer[46]; end
if(wrong_cnt[47] > check_cnt[47]) begin update_buffer[47] <= ~tx_buffer[47]; end else begin update_buffer[47] <= tx_buffer[47]; end
if(wrong_cnt[48] > check_cnt[48]) begin update_buffer[48] <= ~tx_buffer[48]; end else begin update_buffer[48] <= tx_buffer[48]; end
if(wrong_cnt[49] > check_cnt[49]) begin update_buffer[49] <= ~tx_buffer[49]; end else begin update_buffer[49] <= tx_buffer[49]; end
if(wrong_cnt[50] > check_cnt[50]) begin update_buffer[50] <= ~tx_buffer[50]; end else begin update_buffer[50] <= tx_buffer[50]; end
if(wrong_cnt[51] > check_cnt[51]) begin update_buffer[51] <= ~tx_buffer[51]; end else begin update_buffer[51] <= tx_buffer[51]; end
if(wrong_cnt[52] > check_cnt[52]) begin update_buffer[52] <= ~tx_buffer[52]; end else begin update_buffer[52] <= tx_buffer[52]; end
if(wrong_cnt[53] > check_cnt[53]) begin update_buffer[53] <= ~tx_buffer[53]; end else begin update_buffer[53] <= tx_buffer[53]; end
if(wrong_cnt[54] > check_cnt[54]) begin update_buffer[54] <= ~tx_buffer[54]; end else begin update_buffer[54] <= tx_buffer[54]; end
if(wrong_cnt[55] > check_cnt[55]) begin update_buffer[55] <= ~tx_buffer[55]; end else begin update_buffer[55] <= tx_buffer[55]; end
if(wrong_cnt[56] > check_cnt[56]) begin update_buffer[56] <= ~tx_buffer[56]; end else begin update_buffer[56] <= tx_buffer[56]; end
if(wrong_cnt[57] > check_cnt[57]) begin update_buffer[57] <= ~tx_buffer[57]; end else begin update_buffer[57] <= tx_buffer[57]; end
if(wrong_cnt[58] > check_cnt[58]) begin update_buffer[58] <= ~tx_buffer[58]; end else begin update_buffer[58] <= tx_buffer[58]; end
if(wrong_cnt[59] > check_cnt[59]) begin update_buffer[59] <= ~tx_buffer[59]; end else begin update_buffer[59] <= tx_buffer[59]; end
if(wrong_cnt[60] > check_cnt[60]) begin update_buffer[60] <= ~tx_buffer[60]; end else begin update_buffer[60] <= tx_buffer[60]; end
if(wrong_cnt[61] > check_cnt[61]) begin update_buffer[61] <= ~tx_buffer[61]; end else begin update_buffer[61] <= tx_buffer[61]; end
if(wrong_cnt[62] > check_cnt[62]) begin update_buffer[62] <= ~tx_buffer[62]; end else begin update_buffer[62] <= tx_buffer[62]; end
if(wrong_cnt[63] > check_cnt[63]) begin update_buffer[63] <= ~tx_buffer[63]; end else begin update_buffer[63] <= tx_buffer[63]; end
if(wrong_cnt[64] > check_cnt[64]) begin update_buffer[64] <= ~tx_buffer[64]; end else begin update_buffer[64] <= tx_buffer[64]; end
if(wrong_cnt[65] > check_cnt[65]) begin update_buffer[65] <= ~tx_buffer[65]; end else begin update_buffer[65] <= tx_buffer[65]; end
if(wrong_cnt[66] > check_cnt[66]) begin update_buffer[66] <= ~tx_buffer[66]; end else begin update_buffer[66] <= tx_buffer[66]; end
if(wrong_cnt[67] > check_cnt[67]) begin update_buffer[67] <= ~tx_buffer[67]; end else begin update_buffer[67] <= tx_buffer[67]; end
if(wrong_cnt[68] > check_cnt[68]) begin update_buffer[68] <= ~tx_buffer[68]; end else begin update_buffer[68] <= tx_buffer[68]; end
if(wrong_cnt[69] > check_cnt[69]) begin update_buffer[69] <= ~tx_buffer[69]; end else begin update_buffer[69] <= tx_buffer[69]; end
if(wrong_cnt[70] > check_cnt[70]) begin update_buffer[70] <= ~tx_buffer[70]; end else begin update_buffer[70] <= tx_buffer[70]; end
if(wrong_cnt[71] > check_cnt[71]) begin update_buffer[71] <= ~tx_buffer[71]; end else begin update_buffer[71] <= tx_buffer[71]; end
if(wrong_cnt[72] > check_cnt[72]) begin update_buffer[72] <= ~tx_buffer[72]; end else begin update_buffer[72] <= tx_buffer[72]; end
if(wrong_cnt[73] > check_cnt[73]) begin update_buffer[73] <= ~tx_buffer[73]; end else begin update_buffer[73] <= tx_buffer[73]; end
if(wrong_cnt[74] > check_cnt[74]) begin update_buffer[74] <= ~tx_buffer[74]; end else begin update_buffer[74] <= tx_buffer[74]; end
if(wrong_cnt[75] > check_cnt[75]) begin update_buffer[75] <= ~tx_buffer[75]; end else begin update_buffer[75] <= tx_buffer[75]; end
if(wrong_cnt[76] > check_cnt[76]) begin update_buffer[76] <= ~tx_buffer[76]; end else begin update_buffer[76] <= tx_buffer[76]; end
if(wrong_cnt[77] > check_cnt[77]) begin update_buffer[77] <= ~tx_buffer[77]; end else begin update_buffer[77] <= tx_buffer[77]; end
if(wrong_cnt[78] > check_cnt[78]) begin update_buffer[78] <= ~tx_buffer[78]; end else begin update_buffer[78] <= tx_buffer[78]; end
if(wrong_cnt[79] > check_cnt[79]) begin update_buffer[79] <= ~tx_buffer[79]; end else begin update_buffer[79] <= tx_buffer[79]; end
if(wrong_cnt[80] > check_cnt[80]) begin update_buffer[80] <= ~tx_buffer[80]; end else begin update_buffer[80] <= tx_buffer[80]; end
if(wrong_cnt[81] > check_cnt[81]) begin update_buffer[81] <= ~tx_buffer[81]; end else begin update_buffer[81] <= tx_buffer[81]; end
if(wrong_cnt[82] > check_cnt[82]) begin update_buffer[82] <= ~tx_buffer[82]; end else begin update_buffer[82] <= tx_buffer[82]; end
if(wrong_cnt[83] > check_cnt[83]) begin update_buffer[83] <= ~tx_buffer[83]; end else begin update_buffer[83] <= tx_buffer[83]; end
if(wrong_cnt[84] > check_cnt[84]) begin update_buffer[84] <= ~tx_buffer[84]; end else begin update_buffer[84] <= tx_buffer[84]; end
if(wrong_cnt[85] > check_cnt[85]) begin update_buffer[85] <= ~tx_buffer[85]; end else begin update_buffer[85] <= tx_buffer[85]; end
if(wrong_cnt[86] > check_cnt[86]) begin update_buffer[86] <= ~tx_buffer[86]; end else begin update_buffer[86] <= tx_buffer[86]; end
if(wrong_cnt[87] > check_cnt[87]) begin update_buffer[87] <= ~tx_buffer[87]; end else begin update_buffer[87] <= tx_buffer[87]; end
if(wrong_cnt[88] > check_cnt[88]) begin update_buffer[88] <= ~tx_buffer[88]; end else begin update_buffer[88] <= tx_buffer[88]; end
if(wrong_cnt[89] > check_cnt[89]) begin update_buffer[89] <= ~tx_buffer[89]; end else begin update_buffer[89] <= tx_buffer[89]; end
if(wrong_cnt[90] > check_cnt[90]) begin update_buffer[90] <= ~tx_buffer[90]; end else begin update_buffer[90] <= tx_buffer[90]; end
if(wrong_cnt[91] > check_cnt[91]) begin update_buffer[91] <= ~tx_buffer[91]; end else begin update_buffer[91] <= tx_buffer[91]; end
if(wrong_cnt[92] > check_cnt[92]) begin update_buffer[92] <= ~tx_buffer[92]; end else begin update_buffer[92] <= tx_buffer[92]; end
if(wrong_cnt[93] > check_cnt[93]) begin update_buffer[93] <= ~tx_buffer[93]; end else begin update_buffer[93] <= tx_buffer[93]; end
if(wrong_cnt[94] > check_cnt[94]) begin update_buffer[94] <= ~tx_buffer[94]; end else begin update_buffer[94] <= tx_buffer[94]; end
if(wrong_cnt[95] > check_cnt[95]) begin update_buffer[95] <= ~tx_buffer[95]; end else begin update_buffer[95] <= tx_buffer[95]; end
if(wrong_cnt[96] > check_cnt[96]) begin update_buffer[96] <= ~tx_buffer[96]; end else begin update_buffer[96] <= tx_buffer[96]; end
if(wrong_cnt[97] > check_cnt[97]) begin update_buffer[97] <= ~tx_buffer[97]; end else begin update_buffer[97] <= tx_buffer[97]; end
if(wrong_cnt[98] > check_cnt[98]) begin update_buffer[98] <= ~tx_buffer[98]; end else begin update_buffer[98] <= tx_buffer[98]; end
if(wrong_cnt[99] > check_cnt[99]) begin update_buffer[99] <= ~tx_buffer[99]; end else begin update_buffer[99] <= tx_buffer[99]; end
if(wrong_cnt[100] > check_cnt[100]) begin update_buffer[100] <= ~tx_buffer[100]; end else begin update_buffer[100] <= tx_buffer[100]; end
if(wrong_cnt[101] > check_cnt[101]) begin update_buffer[101] <= ~tx_buffer[101]; end else begin update_buffer[101] <= tx_buffer[101]; end
if(wrong_cnt[102] > check_cnt[102]) begin update_buffer[102] <= ~tx_buffer[102]; end else begin update_buffer[102] <= tx_buffer[102]; end
if(wrong_cnt[103] > check_cnt[103]) begin update_buffer[103] <= ~tx_buffer[103]; end else begin update_buffer[103] <= tx_buffer[103]; end
if(wrong_cnt[104] > check_cnt[104]) begin update_buffer[104] <= ~tx_buffer[104]; end else begin update_buffer[104] <= tx_buffer[104]; end
if(wrong_cnt[105] > check_cnt[105]) begin update_buffer[105] <= ~tx_buffer[105]; end else begin update_buffer[105] <= tx_buffer[105]; end
if(wrong_cnt[106] > check_cnt[106]) begin update_buffer[106] <= ~tx_buffer[106]; end else begin update_buffer[106] <= tx_buffer[106]; end
if(wrong_cnt[107] > check_cnt[107]) begin update_buffer[107] <= ~tx_buffer[107]; end else begin update_buffer[107] <= tx_buffer[107]; end
if(wrong_cnt[108] > check_cnt[108]) begin update_buffer[108] <= ~tx_buffer[108]; end else begin update_buffer[108] <= tx_buffer[108]; end
if(wrong_cnt[109] > check_cnt[109]) begin update_buffer[109] <= ~tx_buffer[109]; end else begin update_buffer[109] <= tx_buffer[109]; end
if(wrong_cnt[110] > check_cnt[110]) begin update_buffer[110] <= ~tx_buffer[110]; end else begin update_buffer[110] <= tx_buffer[110]; end
if(wrong_cnt[111] > check_cnt[111]) begin update_buffer[111] <= ~tx_buffer[111]; end else begin update_buffer[111] <= tx_buffer[111]; end
if(wrong_cnt[112] > check_cnt[112]) begin update_buffer[112] <= ~tx_buffer[112]; end else begin update_buffer[112] <= tx_buffer[112]; end
if(wrong_cnt[113] > check_cnt[113]) begin update_buffer[113] <= ~tx_buffer[113]; end else begin update_buffer[113] <= tx_buffer[113]; end
if(wrong_cnt[114] > check_cnt[114]) begin update_buffer[114] <= ~tx_buffer[114]; end else begin update_buffer[114] <= tx_buffer[114]; end
if(wrong_cnt[115] > check_cnt[115]) begin update_buffer[115] <= ~tx_buffer[115]; end else begin update_buffer[115] <= tx_buffer[115]; end
if(wrong_cnt[116] > check_cnt[116]) begin update_buffer[116] <= ~tx_buffer[116]; end else begin update_buffer[116] <= tx_buffer[116]; end
if(wrong_cnt[117] > check_cnt[117]) begin update_buffer[117] <= ~tx_buffer[117]; end else begin update_buffer[117] <= tx_buffer[117]; end
if(wrong_cnt[118] > check_cnt[118]) begin update_buffer[118] <= ~tx_buffer[118]; end else begin update_buffer[118] <= tx_buffer[118]; end
if(wrong_cnt[119] > check_cnt[119]) begin update_buffer[119] <= ~tx_buffer[119]; end else begin update_buffer[119] <= tx_buffer[119]; end
if(wrong_cnt[120] > check_cnt[120]) begin update_buffer[120] <= ~tx_buffer[120]; end else begin update_buffer[120] <= tx_buffer[120]; end
if(wrong_cnt[121] > check_cnt[121]) begin update_buffer[121] <= ~tx_buffer[121]; end else begin update_buffer[121] <= tx_buffer[121]; end
if(wrong_cnt[122] > check_cnt[122]) begin update_buffer[122] <= ~tx_buffer[122]; end else begin update_buffer[122] <= tx_buffer[122]; end
if(wrong_cnt[123] > check_cnt[123]) begin update_buffer[123] <= ~tx_buffer[123]; end else begin update_buffer[123] <= tx_buffer[123]; end
if(wrong_cnt[124] > check_cnt[124]) begin update_buffer[124] <= ~tx_buffer[124]; end else begin update_buffer[124] <= tx_buffer[124]; end
if(wrong_cnt[125] > check_cnt[125]) begin update_buffer[125] <= ~tx_buffer[125]; end else begin update_buffer[125] <= tx_buffer[125]; end
if(wrong_cnt[126] > check_cnt[126]) begin update_buffer[126] <= ~tx_buffer[126]; end else begin update_buffer[126] <= tx_buffer[126]; end
if(wrong_cnt[127] > check_cnt[127]) begin update_buffer[127] <= ~tx_buffer[127]; end else begin update_buffer[127] <= tx_buffer[127]; end
if(wrong_cnt[128] > check_cnt[128]) begin update_buffer[128] <= ~tx_buffer[128]; end else begin update_buffer[128] <= tx_buffer[128]; end
if(wrong_cnt[129] > check_cnt[129]) begin update_buffer[129] <= ~tx_buffer[129]; end else begin update_buffer[129] <= tx_buffer[129]; end
if(wrong_cnt[130] > check_cnt[130]) begin update_buffer[130] <= ~tx_buffer[130]; end else begin update_buffer[130] <= tx_buffer[130]; end
if(wrong_cnt[131] > check_cnt[131]) begin update_buffer[131] <= ~tx_buffer[131]; end else begin update_buffer[131] <= tx_buffer[131]; end
if(wrong_cnt[132] > check_cnt[132]) begin update_buffer[132] <= ~tx_buffer[132]; end else begin update_buffer[132] <= tx_buffer[132]; end
if(wrong_cnt[133] > check_cnt[133]) begin update_buffer[133] <= ~tx_buffer[133]; end else begin update_buffer[133] <= tx_buffer[133]; end
if(wrong_cnt[134] > check_cnt[134]) begin update_buffer[134] <= ~tx_buffer[134]; end else begin update_buffer[134] <= tx_buffer[134]; end
if(wrong_cnt[135] > check_cnt[135]) begin update_buffer[135] <= ~tx_buffer[135]; end else begin update_buffer[135] <= tx_buffer[135]; end
if(wrong_cnt[136] > check_cnt[136]) begin update_buffer[136] <= ~tx_buffer[136]; end else begin update_buffer[136] <= tx_buffer[136]; end
if(wrong_cnt[137] > check_cnt[137]) begin update_buffer[137] <= ~tx_buffer[137]; end else begin update_buffer[137] <= tx_buffer[137]; end
if(wrong_cnt[138] > check_cnt[138]) begin update_buffer[138] <= ~tx_buffer[138]; end else begin update_buffer[138] <= tx_buffer[138]; end
if(wrong_cnt[139] > check_cnt[139]) begin update_buffer[139] <= ~tx_buffer[139]; end else begin update_buffer[139] <= tx_buffer[139]; end
if(wrong_cnt[140] > check_cnt[140]) begin update_buffer[140] <= ~tx_buffer[140]; end else begin update_buffer[140] <= tx_buffer[140]; end
if(wrong_cnt[141] > check_cnt[141]) begin update_buffer[141] <= ~tx_buffer[141]; end else begin update_buffer[141] <= tx_buffer[141]; end
if(wrong_cnt[142] > check_cnt[142]) begin update_buffer[142] <= ~tx_buffer[142]; end else begin update_buffer[142] <= tx_buffer[142]; end
if(wrong_cnt[143] > check_cnt[143]) begin update_buffer[143] <= ~tx_buffer[143]; end else begin update_buffer[143] <= tx_buffer[143]; end
if(wrong_cnt[144] > check_cnt[144]) begin update_buffer[144] <= ~tx_buffer[144]; end else begin update_buffer[144] <= tx_buffer[144]; end
if(wrong_cnt[145] > check_cnt[145]) begin update_buffer[145] <= ~tx_buffer[145]; end else begin update_buffer[145] <= tx_buffer[145]; end
if(wrong_cnt[146] > check_cnt[146]) begin update_buffer[146] <= ~tx_buffer[146]; end else begin update_buffer[146] <= tx_buffer[146]; end
if(wrong_cnt[147] > check_cnt[147]) begin update_buffer[147] <= ~tx_buffer[147]; end else begin update_buffer[147] <= tx_buffer[147]; end
if(wrong_cnt[148] > check_cnt[148]) begin update_buffer[148] <= ~tx_buffer[148]; end else begin update_buffer[148] <= tx_buffer[148]; end
if(wrong_cnt[149] > check_cnt[149]) begin update_buffer[149] <= ~tx_buffer[149]; end else begin update_buffer[149] <= tx_buffer[149]; end
if(wrong_cnt[150] > check_cnt[150]) begin update_buffer[150] <= ~tx_buffer[150]; end else begin update_buffer[150] <= tx_buffer[150]; end
if(wrong_cnt[151] > check_cnt[151]) begin update_buffer[151] <= ~tx_buffer[151]; end else begin update_buffer[151] <= tx_buffer[151]; end
if(wrong_cnt[152] > check_cnt[152]) begin update_buffer[152] <= ~tx_buffer[152]; end else begin update_buffer[152] <= tx_buffer[152]; end
if(wrong_cnt[153] > check_cnt[153]) begin update_buffer[153] <= ~tx_buffer[153]; end else begin update_buffer[153] <= tx_buffer[153]; end
if(wrong_cnt[154] > check_cnt[154]) begin update_buffer[154] <= ~tx_buffer[154]; end else begin update_buffer[154] <= tx_buffer[154]; end
if(wrong_cnt[155] > check_cnt[155]) begin update_buffer[155] <= ~tx_buffer[155]; end else begin update_buffer[155] <= tx_buffer[155]; end
if(wrong_cnt[156] > check_cnt[156]) begin update_buffer[156] <= ~tx_buffer[156]; end else begin update_buffer[156] <= tx_buffer[156]; end
if(wrong_cnt[157] > check_cnt[157]) begin update_buffer[157] <= ~tx_buffer[157]; end else begin update_buffer[157] <= tx_buffer[157]; end
if(wrong_cnt[158] > check_cnt[158]) begin update_buffer[158] <= ~tx_buffer[158]; end else begin update_buffer[158] <= tx_buffer[158]; end
if(wrong_cnt[159] > check_cnt[159]) begin update_buffer[159] <= ~tx_buffer[159]; end else begin update_buffer[159] <= tx_buffer[159]; end
if(wrong_cnt[160] > check_cnt[160]) begin update_buffer[160] <= ~tx_buffer[160]; end else begin update_buffer[160] <= tx_buffer[160]; end
if(wrong_cnt[161] > check_cnt[161]) begin update_buffer[161] <= ~tx_buffer[161]; end else begin update_buffer[161] <= tx_buffer[161]; end
if(wrong_cnt[162] > check_cnt[162]) begin update_buffer[162] <= ~tx_buffer[162]; end else begin update_buffer[162] <= tx_buffer[162]; end
if(wrong_cnt[163] > check_cnt[163]) begin update_buffer[163] <= ~tx_buffer[163]; end else begin update_buffer[163] <= tx_buffer[163]; end
if(wrong_cnt[164] > check_cnt[164]) begin update_buffer[164] <= ~tx_buffer[164]; end else begin update_buffer[164] <= tx_buffer[164]; end
if(wrong_cnt[165] > check_cnt[165]) begin update_buffer[165] <= ~tx_buffer[165]; end else begin update_buffer[165] <= tx_buffer[165]; end
if(wrong_cnt[166] > check_cnt[166]) begin update_buffer[166] <= ~tx_buffer[166]; end else begin update_buffer[166] <= tx_buffer[166]; end
if(wrong_cnt[167] > check_cnt[167]) begin update_buffer[167] <= ~tx_buffer[167]; end else begin update_buffer[167] <= tx_buffer[167]; end
if(wrong_cnt[168] > check_cnt[168]) begin update_buffer[168] <= ~tx_buffer[168]; end else begin update_buffer[168] <= tx_buffer[168]; end
if(wrong_cnt[169] > check_cnt[169]) begin update_buffer[169] <= ~tx_buffer[169]; end else begin update_buffer[169] <= tx_buffer[169]; end
if(wrong_cnt[170] > check_cnt[170]) begin update_buffer[170] <= ~tx_buffer[170]; end else begin update_buffer[170] <= tx_buffer[170]; end
if(wrong_cnt[171] > check_cnt[171]) begin update_buffer[171] <= ~tx_buffer[171]; end else begin update_buffer[171] <= tx_buffer[171]; end
if(wrong_cnt[172] > check_cnt[172]) begin update_buffer[172] <= ~tx_buffer[172]; end else begin update_buffer[172] <= tx_buffer[172]; end
if(wrong_cnt[173] > check_cnt[173]) begin update_buffer[173] <= ~tx_buffer[173]; end else begin update_buffer[173] <= tx_buffer[173]; end
if(wrong_cnt[174] > check_cnt[174]) begin update_buffer[174] <= ~tx_buffer[174]; end else begin update_buffer[174] <= tx_buffer[174]; end
if(wrong_cnt[175] > check_cnt[175]) begin update_buffer[175] <= ~tx_buffer[175]; end else begin update_buffer[175] <= tx_buffer[175]; end
if(wrong_cnt[176] > check_cnt[176]) begin update_buffer[176] <= ~tx_buffer[176]; end else begin update_buffer[176] <= tx_buffer[176]; end
if(wrong_cnt[177] > check_cnt[177]) begin update_buffer[177] <= ~tx_buffer[177]; end else begin update_buffer[177] <= tx_buffer[177]; end
if(wrong_cnt[178] > check_cnt[178]) begin update_buffer[178] <= ~tx_buffer[178]; end else begin update_buffer[178] <= tx_buffer[178]; end
if(wrong_cnt[179] > check_cnt[179]) begin update_buffer[179] <= ~tx_buffer[179]; end else begin update_buffer[179] <= tx_buffer[179]; end
if(wrong_cnt[180] > check_cnt[180]) begin update_buffer[180] <= ~tx_buffer[180]; end else begin update_buffer[180] <= tx_buffer[180]; end
if(wrong_cnt[181] > check_cnt[181]) begin update_buffer[181] <= ~tx_buffer[181]; end else begin update_buffer[181] <= tx_buffer[181]; end
if(wrong_cnt[182] > check_cnt[182]) begin update_buffer[182] <= ~tx_buffer[182]; end else begin update_buffer[182] <= tx_buffer[182]; end
if(wrong_cnt[183] > check_cnt[183]) begin update_buffer[183] <= ~tx_buffer[183]; end else begin update_buffer[183] <= tx_buffer[183]; end
if(wrong_cnt[184] > check_cnt[184]) begin update_buffer[184] <= ~tx_buffer[184]; end else begin update_buffer[184] <= tx_buffer[184]; end
if(wrong_cnt[185] > check_cnt[185]) begin update_buffer[185] <= ~tx_buffer[185]; end else begin update_buffer[185] <= tx_buffer[185]; end
if(wrong_cnt[186] > check_cnt[186]) begin update_buffer[186] <= ~tx_buffer[186]; end else begin update_buffer[186] <= tx_buffer[186]; end
if(wrong_cnt[187] > check_cnt[187]) begin update_buffer[187] <= ~tx_buffer[187]; end else begin update_buffer[187] <= tx_buffer[187]; end
if(wrong_cnt[188] > check_cnt[188]) begin update_buffer[188] <= ~tx_buffer[188]; end else begin update_buffer[188] <= tx_buffer[188]; end
if(wrong_cnt[189] > check_cnt[189]) begin update_buffer[189] <= ~tx_buffer[189]; end else begin update_buffer[189] <= tx_buffer[189]; end
if(wrong_cnt[190] > check_cnt[190]) begin update_buffer[190] <= ~tx_buffer[190]; end else begin update_buffer[190] <= tx_buffer[190]; end
if(wrong_cnt[191] > check_cnt[191]) begin update_buffer[191] <= ~tx_buffer[191]; end else begin update_buffer[191] <= tx_buffer[191]; end
if(wrong_cnt[192] > check_cnt[192]) begin update_buffer[192] <= ~tx_buffer[192]; end else begin update_buffer[192] <= tx_buffer[192]; end
if(wrong_cnt[193] > check_cnt[193]) begin update_buffer[193] <= ~tx_buffer[193]; end else begin update_buffer[193] <= tx_buffer[193]; end
if(wrong_cnt[194] > check_cnt[194]) begin update_buffer[194] <= ~tx_buffer[194]; end else begin update_buffer[194] <= tx_buffer[194]; end
if(wrong_cnt[195] > check_cnt[195]) begin update_buffer[195] <= ~tx_buffer[195]; end else begin update_buffer[195] <= tx_buffer[195]; end
if(wrong_cnt[196] > check_cnt[196]) begin update_buffer[196] <= ~tx_buffer[196]; end else begin update_buffer[196] <= tx_buffer[196]; end
if(wrong_cnt[197] > check_cnt[197]) begin update_buffer[197] <= ~tx_buffer[197]; end else begin update_buffer[197] <= tx_buffer[197]; end
if(wrong_cnt[198] > check_cnt[198]) begin update_buffer[198] <= ~tx_buffer[198]; end else begin update_buffer[198] <= tx_buffer[198]; end
if(wrong_cnt[199] > check_cnt[199]) begin update_buffer[199] <= ~tx_buffer[199]; end else begin update_buffer[199] <= tx_buffer[199]; end
if(wrong_cnt[200] > check_cnt[200]) begin update_buffer[200] <= ~tx_buffer[200]; end else begin update_buffer[200] <= tx_buffer[200]; end
if(wrong_cnt[201] > check_cnt[201]) begin update_buffer[201] <= ~tx_buffer[201]; end else begin update_buffer[201] <= tx_buffer[201]; end
if(wrong_cnt[202] > check_cnt[202]) begin update_buffer[202] <= ~tx_buffer[202]; end else begin update_buffer[202] <= tx_buffer[202]; end
if(wrong_cnt[203] > check_cnt[203]) begin update_buffer[203] <= ~tx_buffer[203]; end else begin update_buffer[203] <= tx_buffer[203]; end
if(wrong_cnt[204] > check_cnt[204]) begin update_buffer[204] <= ~tx_buffer[204]; end else begin update_buffer[204] <= tx_buffer[204]; end
if(wrong_cnt[205] > check_cnt[205]) begin update_buffer[205] <= ~tx_buffer[205]; end else begin update_buffer[205] <= tx_buffer[205]; end
if(wrong_cnt[206] > check_cnt[206]) begin update_buffer[206] <= ~tx_buffer[206]; end else begin update_buffer[206] <= tx_buffer[206]; end
if(wrong_cnt[207] > check_cnt[207]) begin update_buffer[207] <= ~tx_buffer[207]; end else begin update_buffer[207] <= tx_buffer[207]; end
if(wrong_cnt[208] > check_cnt[208]) begin update_buffer[208] <= ~tx_buffer[208]; end else begin update_buffer[208] <= tx_buffer[208]; end
if(wrong_cnt[209] > check_cnt[209]) begin update_buffer[209] <= ~tx_buffer[209]; end else begin update_buffer[209] <= tx_buffer[209]; end
if(wrong_cnt[210] > check_cnt[210]) begin update_buffer[210] <= ~tx_buffer[210]; end else begin update_buffer[210] <= tx_buffer[210]; end
if(wrong_cnt[211] > check_cnt[211]) begin update_buffer[211] <= ~tx_buffer[211]; end else begin update_buffer[211] <= tx_buffer[211]; end
if(wrong_cnt[212] > check_cnt[212]) begin update_buffer[212] <= ~tx_buffer[212]; end else begin update_buffer[212] <= tx_buffer[212]; end
if(wrong_cnt[213] > check_cnt[213]) begin update_buffer[213] <= ~tx_buffer[213]; end else begin update_buffer[213] <= tx_buffer[213]; end
if(wrong_cnt[214] > check_cnt[214]) begin update_buffer[214] <= ~tx_buffer[214]; end else begin update_buffer[214] <= tx_buffer[214]; end
if(wrong_cnt[215] > check_cnt[215]) begin update_buffer[215] <= ~tx_buffer[215]; end else begin update_buffer[215] <= tx_buffer[215]; end
if(wrong_cnt[216] > check_cnt[216]) begin update_buffer[216] <= ~tx_buffer[216]; end else begin update_buffer[216] <= tx_buffer[216]; end
if(wrong_cnt[217] > check_cnt[217]) begin update_buffer[217] <= ~tx_buffer[217]; end else begin update_buffer[217] <= tx_buffer[217]; end
if(wrong_cnt[218] > check_cnt[218]) begin update_buffer[218] <= ~tx_buffer[218]; end else begin update_buffer[218] <= tx_buffer[218]; end
if(wrong_cnt[219] > check_cnt[219]) begin update_buffer[219] <= ~tx_buffer[219]; end else begin update_buffer[219] <= tx_buffer[219]; end
if(wrong_cnt[220] > check_cnt[220]) begin update_buffer[220] <= ~tx_buffer[220]; end else begin update_buffer[220] <= tx_buffer[220]; end
if(wrong_cnt[221] > check_cnt[221]) begin update_buffer[221] <= ~tx_buffer[221]; end else begin update_buffer[221] <= tx_buffer[221]; end
if(wrong_cnt[222] > check_cnt[222]) begin update_buffer[222] <= ~tx_buffer[222]; end else begin update_buffer[222] <= tx_buffer[222]; end
if(wrong_cnt[223] > check_cnt[223]) begin update_buffer[223] <= ~tx_buffer[223]; end else begin update_buffer[223] <= tx_buffer[223]; end
if(wrong_cnt[224] > check_cnt[224]) begin update_buffer[224] <= ~tx_buffer[224]; end else begin update_buffer[224] <= tx_buffer[224]; end
if(wrong_cnt[225] > check_cnt[225]) begin update_buffer[225] <= ~tx_buffer[225]; end else begin update_buffer[225] <= tx_buffer[225]; end
if(wrong_cnt[226] > check_cnt[226]) begin update_buffer[226] <= ~tx_buffer[226]; end else begin update_buffer[226] <= tx_buffer[226]; end
if(wrong_cnt[227] > check_cnt[227]) begin update_buffer[227] <= ~tx_buffer[227]; end else begin update_buffer[227] <= tx_buffer[227]; end
if(wrong_cnt[228] > check_cnt[228]) begin update_buffer[228] <= ~tx_buffer[228]; end else begin update_buffer[228] <= tx_buffer[228]; end
if(wrong_cnt[229] > check_cnt[229]) begin update_buffer[229] <= ~tx_buffer[229]; end else begin update_buffer[229] <= tx_buffer[229]; end
if(wrong_cnt[230] > check_cnt[230]) begin update_buffer[230] <= ~tx_buffer[230]; end else begin update_buffer[230] <= tx_buffer[230]; end
if(wrong_cnt[231] > check_cnt[231]) begin update_buffer[231] <= ~tx_buffer[231]; end else begin update_buffer[231] <= tx_buffer[231]; end
if(wrong_cnt[232] > check_cnt[232]) begin update_buffer[232] <= ~tx_buffer[232]; end else begin update_buffer[232] <= tx_buffer[232]; end
if(wrong_cnt[233] > check_cnt[233]) begin update_buffer[233] <= ~tx_buffer[233]; end else begin update_buffer[233] <= tx_buffer[233]; end
if(wrong_cnt[234] > check_cnt[234]) begin update_buffer[234] <= ~tx_buffer[234]; end else begin update_buffer[234] <= tx_buffer[234]; end
if(wrong_cnt[235] > check_cnt[235]) begin update_buffer[235] <= ~tx_buffer[235]; end else begin update_buffer[235] <= tx_buffer[235]; end
if(wrong_cnt[236] > check_cnt[236]) begin update_buffer[236] <= ~tx_buffer[236]; end else begin update_buffer[236] <= tx_buffer[236]; end
if(wrong_cnt[237] > check_cnt[237]) begin update_buffer[237] <= ~tx_buffer[237]; end else begin update_buffer[237] <= tx_buffer[237]; end
if(wrong_cnt[238] > check_cnt[238]) begin update_buffer[238] <= ~tx_buffer[238]; end else begin update_buffer[238] <= tx_buffer[238]; end
if(wrong_cnt[239] > check_cnt[239]) begin update_buffer[239] <= ~tx_buffer[239]; end else begin update_buffer[239] <= tx_buffer[239]; end
if(wrong_cnt[240] > check_cnt[240]) begin update_buffer[240] <= ~tx_buffer[240]; end else begin update_buffer[240] <= tx_buffer[240]; end
if(wrong_cnt[241] > check_cnt[241]) begin update_buffer[241] <= ~tx_buffer[241]; end else begin update_buffer[241] <= tx_buffer[241]; end
if(wrong_cnt[242] > check_cnt[242]) begin update_buffer[242] <= ~tx_buffer[242]; end else begin update_buffer[242] <= tx_buffer[242]; end
if(wrong_cnt[243] > check_cnt[243]) begin update_buffer[243] <= ~tx_buffer[243]; end else begin update_buffer[243] <= tx_buffer[243]; end
if(wrong_cnt[244] > check_cnt[244]) begin update_buffer[244] <= ~tx_buffer[244]; end else begin update_buffer[244] <= tx_buffer[244]; end
if(wrong_cnt[245] > check_cnt[245]) begin update_buffer[245] <= ~tx_buffer[245]; end else begin update_buffer[245] <= tx_buffer[245]; end
if(wrong_cnt[246] > check_cnt[246]) begin update_buffer[246] <= ~tx_buffer[246]; end else begin update_buffer[246] <= tx_buffer[246]; end
if(wrong_cnt[247] > check_cnt[247]) begin update_buffer[247] <= ~tx_buffer[247]; end else begin update_buffer[247] <= tx_buffer[247]; end
if(wrong_cnt[248] > check_cnt[248]) begin update_buffer[248] <= ~tx_buffer[248]; end else begin update_buffer[248] <= tx_buffer[248]; end
if(wrong_cnt[249] > check_cnt[249]) begin update_buffer[249] <= ~tx_buffer[249]; end else begin update_buffer[249] <= tx_buffer[249]; end
if(wrong_cnt[250] > check_cnt[250]) begin update_buffer[250] <= ~tx_buffer[250]; end else begin update_buffer[250] <= tx_buffer[250]; end
if(wrong_cnt[251] > check_cnt[251]) begin update_buffer[251] <= ~tx_buffer[251]; end else begin update_buffer[251] <= tx_buffer[251]; end
if(wrong_cnt[252] > check_cnt[252]) begin update_buffer[252] <= ~tx_buffer[252]; end else begin update_buffer[252] <= tx_buffer[252]; end
if(wrong_cnt[253] > check_cnt[253]) begin update_buffer[253] <= ~tx_buffer[253]; end else begin update_buffer[253] <= tx_buffer[253]; end
if(wrong_cnt[254] > check_cnt[254]) begin update_buffer[254] <= ~tx_buffer[254]; end else begin update_buffer[254] <= tx_buffer[254]; end
if(wrong_cnt[255] > check_cnt[255]) begin update_buffer[255] <= ~tx_buffer[255]; end else begin update_buffer[255] <= tx_buffer[255]; end

state <= update;

end


update: begin
tx_buffer <= update_buffer;
iter_cnt <= iter_cnt + 1'b1;
if(iter_cnt >= iteration-1) begin
    state <= decode;
end
else begin
    state <= getin;
end

end


decode: begin
valid_flag <= 1'b1;
deout_reg <= tx_buffer;
free_flag <= 1'b1;
iter_cnt <= 'd0;
iter_flag <= 1'b0;
state <= getin;

end

default: state <= init;

endcase


end //the end of biggest if
end //the end of always



endmodule

