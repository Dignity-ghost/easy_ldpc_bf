module add_2.v(a1, a2, s);
input [1:0] a1, a2;
output wire [2:0] s;

assign s = a1 + a2;

endmodule
