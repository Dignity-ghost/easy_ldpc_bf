module add_8(a1, a2, s);
input [3:0] a1, a2;
output wire [4:0] s;

assign s = a1 + a2;

endmodule
