//File name  :    osmlgd_top.v
//Author     :    xiaocuicui
//Time       :    2022/05/21 14:10:24
//Version    :    V1.0
//Abstract   :        


`timescale 1ns/1ps

module osmlgd_top(clk,rst,work,
                  tx,
                  free, deout, valid);

//Define parameters:
parameter iteration = 10;
parameter rigth_formular = 0;

parameter init = 'd0;
parameter getin = 'd1;
parameter dot = 'd2;
parameter judge = 'd3;
parameter check = 'd4;
parameter compare = 'd5;
parameter update = 'd6;
parameter decode = 'd7;

//Define pins:
input clk;
input rst;
input work;
input [255:0] tx;
output wire free;
output wire [255:0] deout;
output wire valid;

//Define signals:
reg [2:0] state;

reg [255:0] Harray [127:0];
reg [255:0] tx_buffer;
reg [255:0] dotarray [127:0];
reg [127:0] form_array;
reg [7:0] check_cnt [255:0];
reg [7:0] wrong_cnt [255:0];
reg [255:0] update_buffer;
reg [3:0] iter_cnt;
reg free_flag, valid_flag, iter_flag;
reg [255:0] deout_reg;

assign free = free_flag;
assign valid = valid_flag;
assign deout = deout_reg;

//Instance

wire [8:0] row_sum_0, row_sum_1, row_sum_2, row_sum_3, row_sum_4, row_sum_5, row_sum_6, row_sum_7, 
           row_sum_8, row_sum_9, row_sum_10, row_sum_11, row_sum_12, row_sum_13, row_sum_14, row_sum_15, 
           row_sum_16, row_sum_17, row_sum_18, row_sum_19, row_sum_20, row_sum_21, row_sum_22, row_sum_23, 
           row_sum_24, row_sum_25, row_sum_26, row_sum_27, row_sum_28, row_sum_29, row_sum_30, row_sum_31, 
           row_sum_32, row_sum_33, row_sum_34, row_sum_35, row_sum_36, row_sum_37, row_sum_38, row_sum_39, 
           row_sum_40, row_sum_41, row_sum_42, row_sum_43, row_sum_44, row_sum_45, row_sum_46, row_sum_47, 
           row_sum_48, row_sum_49, row_sum_50, row_sum_51, row_sum_52, row_sum_53, row_sum_54, row_sum_55, 
           row_sum_56, row_sum_57, row_sum_58, row_sum_59, row_sum_60, row_sum_61, row_sum_62, row_sum_63, 
           row_sum_64, row_sum_65, row_sum_66, row_sum_67, row_sum_68, row_sum_69, row_sum_70, row_sum_71, 
           row_sum_72, row_sum_73, row_sum_74, row_sum_75, row_sum_76, row_sum_77, row_sum_78, row_sum_79, 
           row_sum_80, row_sum_81, row_sum_82, row_sum_83, row_sum_84, row_sum_85, row_sum_86, row_sum_87, 
           row_sum_88, row_sum_89, row_sum_90, row_sum_91, row_sum_92, row_sum_93, row_sum_94, row_sum_95, 
           row_sum_96, row_sum_97, row_sum_98, row_sum_99, row_sum_100, row_sum_101, row_sum_102, row_sum_103, 
           row_sum_104, row_sum_105, row_sum_106, row_sum_107, row_sum_108, row_sum_109, row_sum_110, row_sum_111, 
           row_sum_112, row_sum_113, row_sum_114, row_sum_115, row_sum_116, row_sum_117, row_sum_118, row_sum_119, 
           row_sum_120, row_sum_121, row_sum_122, row_sum_123, row_sum_124, row_sum_125, row_sum_126, row_sum_127;

wire [127:0] row_sum_lastbit;

assign row_sum_lastbit = {row_sum_127[0], row_sum_126[0], row_sum_125[0], row_sum_124[0], row_sum_123[0], row_sum_122[0], row_sum_121[0], row_sum_120[0], 
                          row_sum_119[0], row_sum_118[0], row_sum_117[0], row_sum_116[0], row_sum_115[0], row_sum_114[0], row_sum_113[0], row_sum_112[0], 
                          row_sum_111[0], row_sum_110[0], row_sum_109[0], row_sum_108[0], row_sum_107[0], row_sum_106[0], row_sum_105[0], row_sum_104[0], 
                          row_sum_103[0], row_sum_102[0], row_sum_101[0], row_sum_100[0], row_sum_99[0], row_sum_98[0], row_sum_97[0], row_sum_96[0], 
                          row_sum_95[0], row_sum_94[0], row_sum_93[0], row_sum_92[0], row_sum_91[0], row_sum_90[0], row_sum_89[0], row_sum_88[0], 
                          row_sum_87[0], row_sum_86[0], row_sum_85[0], row_sum_84[0], row_sum_83[0], row_sum_82[0], row_sum_81[0], row_sum_80[0], 
                          row_sum_79[0], row_sum_78[0], row_sum_77[0], row_sum_76[0], row_sum_75[0], row_sum_74[0], row_sum_73[0], row_sum_72[0], 
                          row_sum_71[0], row_sum_70[0], row_sum_69[0], row_sum_68[0], row_sum_67[0], row_sum_66[0], row_sum_65[0], row_sum_64[0], 
                          row_sum_63[0], row_sum_62[0], row_sum_61[0], row_sum_60[0], row_sum_59[0], row_sum_58[0], row_sum_57[0], row_sum_56[0], 
                          row_sum_55[0], row_sum_54[0], row_sum_53[0], row_sum_52[0], row_sum_51[0], row_sum_50[0], row_sum_49[0], row_sum_48[0], 
                          row_sum_47[0], row_sum_46[0], row_sum_45[0], row_sum_44[0], row_sum_43[0], row_sum_42[0], row_sum_41[0], row_sum_40[0], 
                          row_sum_39[0], row_sum_38[0], row_sum_37[0], row_sum_36[0], row_sum_35[0], row_sum_34[0], row_sum_33[0], row_sum_32[0], 
                          row_sum_31[0], row_sum_30[0], row_sum_29[0], row_sum_28[0], row_sum_27[0], row_sum_26[0], row_sum_25[0], row_sum_24[0], 
                          row_sum_23[0], row_sum_22[0], row_sum_21[0], row_sum_20[0], row_sum_19[0], row_sum_18[0], row_sum_17[0], row_sum_16[0], 
                          row_sum_15[0], row_sum_14[0], row_sum_13[0], row_sum_12[0], row_sum_11[0], row_sum_10[0], row_sum_9[0], row_sum_8[0], 
                          row_sum_7[0], row_sum_6[0], row_sum_5[0], row_sum_4[0], row_sum_3[0], row_sum_2[0], row_sum_1[0], row_sum_0[0]};


bitsadder_256 f_check_0(dotarray[0], row_sum_0);
bitsadder_256 f_check_1(dotarray[1], row_sum_1);
bitsadder_256 f_check_2(dotarray[2], row_sum_2);
bitsadder_256 f_check_3(dotarray[3], row_sum_3);
bitsadder_256 f_check_4(dotarray[4], row_sum_4);
bitsadder_256 f_check_5(dotarray[5], row_sum_5);
bitsadder_256 f_check_6(dotarray[6], row_sum_6);
bitsadder_256 f_check_7(dotarray[7], row_sum_7);
bitsadder_256 f_check_8(dotarray[8], row_sum_8);
bitsadder_256 f_check_9(dotarray[9], row_sum_9);
bitsadder_256 f_check_10(dotarray[10], row_sum_10);
bitsadder_256 f_check_11(dotarray[11], row_sum_11);
bitsadder_256 f_check_12(dotarray[12], row_sum_12);
bitsadder_256 f_check_13(dotarray[13], row_sum_13);
bitsadder_256 f_check_14(dotarray[14], row_sum_14);
bitsadder_256 f_check_15(dotarray[15], row_sum_15);
bitsadder_256 f_check_16(dotarray[16], row_sum_16);
bitsadder_256 f_check_17(dotarray[17], row_sum_17);
bitsadder_256 f_check_18(dotarray[18], row_sum_18);
bitsadder_256 f_check_19(dotarray[19], row_sum_19);
bitsadder_256 f_check_20(dotarray[20], row_sum_20);
bitsadder_256 f_check_21(dotarray[21], row_sum_21);
bitsadder_256 f_check_22(dotarray[22], row_sum_22);
bitsadder_256 f_check_23(dotarray[23], row_sum_23);
bitsadder_256 f_check_24(dotarray[24], row_sum_24);
bitsadder_256 f_check_25(dotarray[25], row_sum_25);
bitsadder_256 f_check_26(dotarray[26], row_sum_26);
bitsadder_256 f_check_27(dotarray[27], row_sum_27);
bitsadder_256 f_check_28(dotarray[28], row_sum_28);
bitsadder_256 f_check_29(dotarray[29], row_sum_29);
bitsadder_256 f_check_30(dotarray[30], row_sum_30);
bitsadder_256 f_check_31(dotarray[31], row_sum_31);
bitsadder_256 f_check_32(dotarray[32], row_sum_32);
bitsadder_256 f_check_33(dotarray[33], row_sum_33);
bitsadder_256 f_check_34(dotarray[34], row_sum_34);
bitsadder_256 f_check_35(dotarray[35], row_sum_35);
bitsadder_256 f_check_36(dotarray[36], row_sum_36);
bitsadder_256 f_check_37(dotarray[37], row_sum_37);
bitsadder_256 f_check_38(dotarray[38], row_sum_38);
bitsadder_256 f_check_39(dotarray[39], row_sum_39);
bitsadder_256 f_check_40(dotarray[40], row_sum_40);
bitsadder_256 f_check_41(dotarray[41], row_sum_41);
bitsadder_256 f_check_42(dotarray[42], row_sum_42);
bitsadder_256 f_check_43(dotarray[43], row_sum_43);
bitsadder_256 f_check_44(dotarray[44], row_sum_44);
bitsadder_256 f_check_45(dotarray[45], row_sum_45);
bitsadder_256 f_check_46(dotarray[46], row_sum_46);
bitsadder_256 f_check_47(dotarray[47], row_sum_47);
bitsadder_256 f_check_48(dotarray[48], row_sum_48);
bitsadder_256 f_check_49(dotarray[49], row_sum_49);
bitsadder_256 f_check_50(dotarray[50], row_sum_50);
bitsadder_256 f_check_51(dotarray[51], row_sum_51);
bitsadder_256 f_check_52(dotarray[52], row_sum_52);
bitsadder_256 f_check_53(dotarray[53], row_sum_53);
bitsadder_256 f_check_54(dotarray[54], row_sum_54);
bitsadder_256 f_check_55(dotarray[55], row_sum_55);
bitsadder_256 f_check_56(dotarray[56], row_sum_56);
bitsadder_256 f_check_57(dotarray[57], row_sum_57);
bitsadder_256 f_check_58(dotarray[58], row_sum_58);
bitsadder_256 f_check_59(dotarray[59], row_sum_59);
bitsadder_256 f_check_60(dotarray[60], row_sum_60);
bitsadder_256 f_check_61(dotarray[61], row_sum_61);
bitsadder_256 f_check_62(dotarray[62], row_sum_62);
bitsadder_256 f_check_63(dotarray[63], row_sum_63);
bitsadder_256 f_check_64(dotarray[64], row_sum_64);
bitsadder_256 f_check_65(dotarray[65], row_sum_65);
bitsadder_256 f_check_66(dotarray[66], row_sum_66);
bitsadder_256 f_check_67(dotarray[67], row_sum_67);
bitsadder_256 f_check_68(dotarray[68], row_sum_68);
bitsadder_256 f_check_69(dotarray[69], row_sum_69);
bitsadder_256 f_check_70(dotarray[70], row_sum_70);
bitsadder_256 f_check_71(dotarray[71], row_sum_71);
bitsadder_256 f_check_72(dotarray[72], row_sum_72);
bitsadder_256 f_check_73(dotarray[73], row_sum_73);
bitsadder_256 f_check_74(dotarray[74], row_sum_74);
bitsadder_256 f_check_75(dotarray[75], row_sum_75);
bitsadder_256 f_check_76(dotarray[76], row_sum_76);
bitsadder_256 f_check_77(dotarray[77], row_sum_77);
bitsadder_256 f_check_78(dotarray[78], row_sum_78);
bitsadder_256 f_check_79(dotarray[79], row_sum_79);
bitsadder_256 f_check_80(dotarray[80], row_sum_80);
bitsadder_256 f_check_81(dotarray[81], row_sum_81);
bitsadder_256 f_check_82(dotarray[82], row_sum_82);
bitsadder_256 f_check_83(dotarray[83], row_sum_83);
bitsadder_256 f_check_84(dotarray[84], row_sum_84);
bitsadder_256 f_check_85(dotarray[85], row_sum_85);
bitsadder_256 f_check_86(dotarray[86], row_sum_86);
bitsadder_256 f_check_87(dotarray[87], row_sum_87);
bitsadder_256 f_check_88(dotarray[88], row_sum_88);
bitsadder_256 f_check_89(dotarray[89], row_sum_89);
bitsadder_256 f_check_90(dotarray[90], row_sum_90);
bitsadder_256 f_check_91(dotarray[91], row_sum_91);
bitsadder_256 f_check_92(dotarray[92], row_sum_92);
bitsadder_256 f_check_93(dotarray[93], row_sum_93);
bitsadder_256 f_check_94(dotarray[94], row_sum_94);
bitsadder_256 f_check_95(dotarray[95], row_sum_95);
bitsadder_256 f_check_96(dotarray[96], row_sum_96);
bitsadder_256 f_check_97(dotarray[97], row_sum_97);
bitsadder_256 f_check_98(dotarray[98], row_sum_98);
bitsadder_256 f_check_99(dotarray[99], row_sum_99);
bitsadder_256 f_check_100(dotarray[100], row_sum_100);
bitsadder_256 f_check_101(dotarray[101], row_sum_101);
bitsadder_256 f_check_102(dotarray[102], row_sum_102);
bitsadder_256 f_check_103(dotarray[103], row_sum_103);
bitsadder_256 f_check_104(dotarray[104], row_sum_104);
bitsadder_256 f_check_105(dotarray[105], row_sum_105);
bitsadder_256 f_check_106(dotarray[106], row_sum_106);
bitsadder_256 f_check_107(dotarray[107], row_sum_107);
bitsadder_256 f_check_108(dotarray[108], row_sum_108);
bitsadder_256 f_check_109(dotarray[109], row_sum_109);
bitsadder_256 f_check_110(dotarray[110], row_sum_110);
bitsadder_256 f_check_111(dotarray[111], row_sum_111);
bitsadder_256 f_check_112(dotarray[112], row_sum_112);
bitsadder_256 f_check_113(dotarray[113], row_sum_113);
bitsadder_256 f_check_114(dotarray[114], row_sum_114);
bitsadder_256 f_check_115(dotarray[115], row_sum_115);
bitsadder_256 f_check_116(dotarray[116], row_sum_116);
bitsadder_256 f_check_117(dotarray[117], row_sum_117);
bitsadder_256 f_check_118(dotarray[118], row_sum_118);
bitsadder_256 f_check_119(dotarray[119], row_sum_119);
bitsadder_256 f_check_120(dotarray[120], row_sum_120);
bitsadder_256 f_check_121(dotarray[121], row_sum_121);
bitsadder_256 f_check_122(dotarray[122], row_sum_122);
bitsadder_256 f_check_123(dotarray[123], row_sum_123);
bitsadder_256 f_check_124(dotarray[124], row_sum_124);
bitsadder_256 f_check_125(dotarray[125], row_sum_125);
bitsadder_256 f_check_126(dotarray[126], row_sum_126);
bitsadder_256 f_check_127(dotarray[127], row_sum_127);


wire [127:0] dot_col_0, dot_col_1, dot_col_2, dot_col_3, dot_col_4, dot_col_5, dot_col_6, dot_col_7, 
             dot_col_8, dot_col_9, dot_col_10, dot_col_11, dot_col_12, dot_col_13, dot_col_14, dot_col_15, 
             dot_col_16, dot_col_17, dot_col_18, dot_col_19, dot_col_20, dot_col_21, dot_col_22, dot_col_23, 
             dot_col_24, dot_col_25, dot_col_26, dot_col_27, dot_col_28, dot_col_29, dot_col_30, dot_col_31, 
             dot_col_32, dot_col_33, dot_col_34, dot_col_35, dot_col_36, dot_col_37, dot_col_38, dot_col_39, 
             dot_col_40, dot_col_41, dot_col_42, dot_col_43, dot_col_44, dot_col_45, dot_col_46, dot_col_47, 
             dot_col_48, dot_col_49, dot_col_50, dot_col_51, dot_col_52, dot_col_53, dot_col_54, dot_col_55, 
             dot_col_56, dot_col_57, dot_col_58, dot_col_59, dot_col_60, dot_col_61, dot_col_62, dot_col_63, 
             dot_col_64, dot_col_65, dot_col_66, dot_col_67, dot_col_68, dot_col_69, dot_col_70, dot_col_71, 
             dot_col_72, dot_col_73, dot_col_74, dot_col_75, dot_col_76, dot_col_77, dot_col_78, dot_col_79, 
             dot_col_80, dot_col_81, dot_col_82, dot_col_83, dot_col_84, dot_col_85, dot_col_86, dot_col_87, 
             dot_col_88, dot_col_89, dot_col_90, dot_col_91, dot_col_92, dot_col_93, dot_col_94, dot_col_95, 
             dot_col_96, dot_col_97, dot_col_98, dot_col_99, dot_col_100, dot_col_101, dot_col_102, dot_col_103, 
             dot_col_104, dot_col_105, dot_col_106, dot_col_107, dot_col_108, dot_col_109, dot_col_110, dot_col_111, 
             dot_col_112, dot_col_113, dot_col_114, dot_col_115, dot_col_116, dot_col_117, dot_col_118, dot_col_119, 
             dot_col_120, dot_col_121, dot_col_122, dot_col_123, dot_col_124, dot_col_125, dot_col_126, dot_col_127, 
             dot_col_128, dot_col_129, dot_col_130, dot_col_131, dot_col_132, dot_col_133, dot_col_134, dot_col_135, 
             dot_col_136, dot_col_137, dot_col_138, dot_col_139, dot_col_140, dot_col_141, dot_col_142, dot_col_143, 
             dot_col_144, dot_col_145, dot_col_146, dot_col_147, dot_col_148, dot_col_149, dot_col_150, dot_col_151, 
             dot_col_152, dot_col_153, dot_col_154, dot_col_155, dot_col_156, dot_col_157, dot_col_158, dot_col_159, 
             dot_col_160, dot_col_161, dot_col_162, dot_col_163, dot_col_164, dot_col_165, dot_col_166, dot_col_167, 
             dot_col_168, dot_col_169, dot_col_170, dot_col_171, dot_col_172, dot_col_173, dot_col_174, dot_col_175, 
             dot_col_176, dot_col_177, dot_col_178, dot_col_179, dot_col_180, dot_col_181, dot_col_182, dot_col_183, 
             dot_col_184, dot_col_185, dot_col_186, dot_col_187, dot_col_188, dot_col_189, dot_col_190, dot_col_191, 
             dot_col_192, dot_col_193, dot_col_194, dot_col_195, dot_col_196, dot_col_197, dot_col_198, dot_col_199, 
             dot_col_200, dot_col_201, dot_col_202, dot_col_203, dot_col_204, dot_col_205, dot_col_206, dot_col_207, 
             dot_col_208, dot_col_209, dot_col_210, dot_col_211, dot_col_212, dot_col_213, dot_col_214, dot_col_215, 
             dot_col_216, dot_col_217, dot_col_218, dot_col_219, dot_col_220, dot_col_221, dot_col_222, dot_col_223, 
             dot_col_224, dot_col_225, dot_col_226, dot_col_227, dot_col_228, dot_col_229, dot_col_230, dot_col_231, 
             dot_col_232, dot_col_233, dot_col_234, dot_col_235, dot_col_236, dot_col_237, dot_col_238, dot_col_239, 
             dot_col_240, dot_col_241, dot_col_242, dot_col_243, dot_col_244, dot_col_245, dot_col_246, dot_col_247, 
             dot_col_248, dot_col_249, dot_col_250, dot_col_251, dot_col_252, dot_col_253, dot_col_254, dot_col_255;

assign dot_col_0 = {dotarray[0][0], dotarray[1][0], dotarray[2][0], dotarray[3][0], dotarray[4][0], dotarray[5][0], dotarray[6][0], dotarray[7][0], dotarray[8][0], dotarray[9][0], dotarray[10][0], dotarray[11][0], dotarray[12][0], dotarray[13][0], dotarray[14][0], dotarray[15][0], dotarray[16][0], dotarray[17][0], dotarray[18][0], dotarray[19][0], dotarray[20][0], dotarray[21][0], dotarray[22][0], dotarray[23][0], dotarray[24][0], dotarray[25][0], dotarray[26][0], dotarray[27][0], dotarray[28][0], dotarray[29][0], dotarray[30][0], dotarray[31][0], dotarray[32][0], dotarray[33][0], dotarray[34][0], dotarray[35][0], dotarray[36][0], dotarray[37][0], dotarray[38][0], dotarray[39][0], dotarray[40][0], dotarray[41][0], dotarray[42][0], dotarray[43][0], dotarray[44][0], dotarray[45][0], dotarray[46][0], dotarray[47][0], dotarray[48][0], dotarray[49][0], dotarray[50][0], dotarray[51][0], dotarray[52][0], dotarray[53][0], dotarray[54][0], dotarray[55][0], dotarray[56][0], dotarray[57][0], dotarray[58][0], dotarray[59][0], dotarray[60][0], dotarray[61][0], dotarray[62][0], dotarray[63][0], dotarray[64][0], dotarray[65][0], dotarray[66][0], dotarray[67][0], dotarray[68][0], dotarray[69][0], dotarray[70][0], dotarray[71][0], dotarray[72][0], dotarray[73][0], dotarray[74][0], dotarray[75][0], dotarray[76][0], dotarray[77][0], dotarray[78][0], dotarray[79][0], dotarray[80][0], dotarray[81][0], dotarray[82][0], dotarray[83][0], dotarray[84][0], dotarray[85][0], dotarray[86][0], dotarray[87][0], dotarray[88][0], dotarray[89][0], dotarray[90][0], dotarray[91][0], dotarray[92][0], dotarray[93][0], dotarray[94][0], dotarray[95][0], dotarray[96][0], dotarray[97][0], dotarray[98][0], dotarray[99][0], dotarray[100][0], dotarray[101][0], dotarray[102][0], dotarray[103][0], dotarray[104][0], dotarray[105][0], dotarray[106][0], dotarray[107][0], dotarray[108][0], dotarray[109][0], dotarray[110][0], dotarray[111][0], dotarray[112][0], dotarray[113][0], dotarray[114][0], dotarray[115][0], dotarray[116][0], dotarray[117][0], dotarray[118][0], dotarray[119][0], dotarray[120][0], dotarray[121][0], dotarray[122][0], dotarray[123][0], dotarray[124][0], dotarray[125][0], dotarray[126][0], dotarray[127][0]};
assign dot_col_1 = {dotarray[0][1], dotarray[1][1], dotarray[2][1], dotarray[3][1], dotarray[4][1], dotarray[5][1], dotarray[6][1], dotarray[7][1], dotarray[8][1], dotarray[9][1], dotarray[10][1], dotarray[11][1], dotarray[12][1], dotarray[13][1], dotarray[14][1], dotarray[15][1], dotarray[16][1], dotarray[17][1], dotarray[18][1], dotarray[19][1], dotarray[20][1], dotarray[21][1], dotarray[22][1], dotarray[23][1], dotarray[24][1], dotarray[25][1], dotarray[26][1], dotarray[27][1], dotarray[28][1], dotarray[29][1], dotarray[30][1], dotarray[31][1], dotarray[32][1], dotarray[33][1], dotarray[34][1], dotarray[35][1], dotarray[36][1], dotarray[37][1], dotarray[38][1], dotarray[39][1], dotarray[40][1], dotarray[41][1], dotarray[42][1], dotarray[43][1], dotarray[44][1], dotarray[45][1], dotarray[46][1], dotarray[47][1], dotarray[48][1], dotarray[49][1], dotarray[50][1], dotarray[51][1], dotarray[52][1], dotarray[53][1], dotarray[54][1], dotarray[55][1], dotarray[56][1], dotarray[57][1], dotarray[58][1], dotarray[59][1], dotarray[60][1], dotarray[61][1], dotarray[62][1], dotarray[63][1], dotarray[64][1], dotarray[65][1], dotarray[66][1], dotarray[67][1], dotarray[68][1], dotarray[69][1], dotarray[70][1], dotarray[71][1], dotarray[72][1], dotarray[73][1], dotarray[74][1], dotarray[75][1], dotarray[76][1], dotarray[77][1], dotarray[78][1], dotarray[79][1], dotarray[80][1], dotarray[81][1], dotarray[82][1], dotarray[83][1], dotarray[84][1], dotarray[85][1], dotarray[86][1], dotarray[87][1], dotarray[88][1], dotarray[89][1], dotarray[90][1], dotarray[91][1], dotarray[92][1], dotarray[93][1], dotarray[94][1], dotarray[95][1], dotarray[96][1], dotarray[97][1], dotarray[98][1], dotarray[99][1], dotarray[100][1], dotarray[101][1], dotarray[102][1], dotarray[103][1], dotarray[104][1], dotarray[105][1], dotarray[106][1], dotarray[107][1], dotarray[108][1], dotarray[109][1], dotarray[110][1], dotarray[111][1], dotarray[112][1], dotarray[113][1], dotarray[114][1], dotarray[115][1], dotarray[116][1], dotarray[117][1], dotarray[118][1], dotarray[119][1], dotarray[120][1], dotarray[121][1], dotarray[122][1], dotarray[123][1], dotarray[124][1], dotarray[125][1], dotarray[126][1], dotarray[127][1]};
assign dot_col_2 = {dotarray[0][2], dotarray[1][2], dotarray[2][2], dotarray[3][2], dotarray[4][2], dotarray[5][2], dotarray[6][2], dotarray[7][2], dotarray[8][2], dotarray[9][2], dotarray[10][2], dotarray[11][2], dotarray[12][2], dotarray[13][2], dotarray[14][2], dotarray[15][2], dotarray[16][2], dotarray[17][2], dotarray[18][2], dotarray[19][2], dotarray[20][2], dotarray[21][2], dotarray[22][2], dotarray[23][2], dotarray[24][2], dotarray[25][2], dotarray[26][2], dotarray[27][2], dotarray[28][2], dotarray[29][2], dotarray[30][2], dotarray[31][2], dotarray[32][2], dotarray[33][2], dotarray[34][2], dotarray[35][2], dotarray[36][2], dotarray[37][2], dotarray[38][2], dotarray[39][2], dotarray[40][2], dotarray[41][2], dotarray[42][2], dotarray[43][2], dotarray[44][2], dotarray[45][2], dotarray[46][2], dotarray[47][2], dotarray[48][2], dotarray[49][2], dotarray[50][2], dotarray[51][2], dotarray[52][2], dotarray[53][2], dotarray[54][2], dotarray[55][2], dotarray[56][2], dotarray[57][2], dotarray[58][2], dotarray[59][2], dotarray[60][2], dotarray[61][2], dotarray[62][2], dotarray[63][2], dotarray[64][2], dotarray[65][2], dotarray[66][2], dotarray[67][2], dotarray[68][2], dotarray[69][2], dotarray[70][2], dotarray[71][2], dotarray[72][2], dotarray[73][2], dotarray[74][2], dotarray[75][2], dotarray[76][2], dotarray[77][2], dotarray[78][2], dotarray[79][2], dotarray[80][2], dotarray[81][2], dotarray[82][2], dotarray[83][2], dotarray[84][2], dotarray[85][2], dotarray[86][2], dotarray[87][2], dotarray[88][2], dotarray[89][2], dotarray[90][2], dotarray[91][2], dotarray[92][2], dotarray[93][2], dotarray[94][2], dotarray[95][2], dotarray[96][2], dotarray[97][2], dotarray[98][2], dotarray[99][2], dotarray[100][2], dotarray[101][2], dotarray[102][2], dotarray[103][2], dotarray[104][2], dotarray[105][2], dotarray[106][2], dotarray[107][2], dotarray[108][2], dotarray[109][2], dotarray[110][2], dotarray[111][2], dotarray[112][2], dotarray[113][2], dotarray[114][2], dotarray[115][2], dotarray[116][2], dotarray[117][2], dotarray[118][2], dotarray[119][2], dotarray[120][2], dotarray[121][2], dotarray[122][2], dotarray[123][2], dotarray[124][2], dotarray[125][2], dotarray[126][2], dotarray[127][2]};
assign dot_col_3 = {dotarray[0][3], dotarray[1][3], dotarray[2][3], dotarray[3][3], dotarray[4][3], dotarray[5][3], dotarray[6][3], dotarray[7][3], dotarray[8][3], dotarray[9][3], dotarray[10][3], dotarray[11][3], dotarray[12][3], dotarray[13][3], dotarray[14][3], dotarray[15][3], dotarray[16][3], dotarray[17][3], dotarray[18][3], dotarray[19][3], dotarray[20][3], dotarray[21][3], dotarray[22][3], dotarray[23][3], dotarray[24][3], dotarray[25][3], dotarray[26][3], dotarray[27][3], dotarray[28][3], dotarray[29][3], dotarray[30][3], dotarray[31][3], dotarray[32][3], dotarray[33][3], dotarray[34][3], dotarray[35][3], dotarray[36][3], dotarray[37][3], dotarray[38][3], dotarray[39][3], dotarray[40][3], dotarray[41][3], dotarray[42][3], dotarray[43][3], dotarray[44][3], dotarray[45][3], dotarray[46][3], dotarray[47][3], dotarray[48][3], dotarray[49][3], dotarray[50][3], dotarray[51][3], dotarray[52][3], dotarray[53][3], dotarray[54][3], dotarray[55][3], dotarray[56][3], dotarray[57][3], dotarray[58][3], dotarray[59][3], dotarray[60][3], dotarray[61][3], dotarray[62][3], dotarray[63][3], dotarray[64][3], dotarray[65][3], dotarray[66][3], dotarray[67][3], dotarray[68][3], dotarray[69][3], dotarray[70][3], dotarray[71][3], dotarray[72][3], dotarray[73][3], dotarray[74][3], dotarray[75][3], dotarray[76][3], dotarray[77][3], dotarray[78][3], dotarray[79][3], dotarray[80][3], dotarray[81][3], dotarray[82][3], dotarray[83][3], dotarray[84][3], dotarray[85][3], dotarray[86][3], dotarray[87][3], dotarray[88][3], dotarray[89][3], dotarray[90][3], dotarray[91][3], dotarray[92][3], dotarray[93][3], dotarray[94][3], dotarray[95][3], dotarray[96][3], dotarray[97][3], dotarray[98][3], dotarray[99][3], dotarray[100][3], dotarray[101][3], dotarray[102][3], dotarray[103][3], dotarray[104][3], dotarray[105][3], dotarray[106][3], dotarray[107][3], dotarray[108][3], dotarray[109][3], dotarray[110][3], dotarray[111][3], dotarray[112][3], dotarray[113][3], dotarray[114][3], dotarray[115][3], dotarray[116][3], dotarray[117][3], dotarray[118][3], dotarray[119][3], dotarray[120][3], dotarray[121][3], dotarray[122][3], dotarray[123][3], dotarray[124][3], dotarray[125][3], dotarray[126][3], dotarray[127][3]};
assign dot_col_4 = {dotarray[0][4], dotarray[1][4], dotarray[2][4], dotarray[3][4], dotarray[4][4], dotarray[5][4], dotarray[6][4], dotarray[7][4], dotarray[8][4], dotarray[9][4], dotarray[10][4], dotarray[11][4], dotarray[12][4], dotarray[13][4], dotarray[14][4], dotarray[15][4], dotarray[16][4], dotarray[17][4], dotarray[18][4], dotarray[19][4], dotarray[20][4], dotarray[21][4], dotarray[22][4], dotarray[23][4], dotarray[24][4], dotarray[25][4], dotarray[26][4], dotarray[27][4], dotarray[28][4], dotarray[29][4], dotarray[30][4], dotarray[31][4], dotarray[32][4], dotarray[33][4], dotarray[34][4], dotarray[35][4], dotarray[36][4], dotarray[37][4], dotarray[38][4], dotarray[39][4], dotarray[40][4], dotarray[41][4], dotarray[42][4], dotarray[43][4], dotarray[44][4], dotarray[45][4], dotarray[46][4], dotarray[47][4], dotarray[48][4], dotarray[49][4], dotarray[50][4], dotarray[51][4], dotarray[52][4], dotarray[53][4], dotarray[54][4], dotarray[55][4], dotarray[56][4], dotarray[57][4], dotarray[58][4], dotarray[59][4], dotarray[60][4], dotarray[61][4], dotarray[62][4], dotarray[63][4], dotarray[64][4], dotarray[65][4], dotarray[66][4], dotarray[67][4], dotarray[68][4], dotarray[69][4], dotarray[70][4], dotarray[71][4], dotarray[72][4], dotarray[73][4], dotarray[74][4], dotarray[75][4], dotarray[76][4], dotarray[77][4], dotarray[78][4], dotarray[79][4], dotarray[80][4], dotarray[81][4], dotarray[82][4], dotarray[83][4], dotarray[84][4], dotarray[85][4], dotarray[86][4], dotarray[87][4], dotarray[88][4], dotarray[89][4], dotarray[90][4], dotarray[91][4], dotarray[92][4], dotarray[93][4], dotarray[94][4], dotarray[95][4], dotarray[96][4], dotarray[97][4], dotarray[98][4], dotarray[99][4], dotarray[100][4], dotarray[101][4], dotarray[102][4], dotarray[103][4], dotarray[104][4], dotarray[105][4], dotarray[106][4], dotarray[107][4], dotarray[108][4], dotarray[109][4], dotarray[110][4], dotarray[111][4], dotarray[112][4], dotarray[113][4], dotarray[114][4], dotarray[115][4], dotarray[116][4], dotarray[117][4], dotarray[118][4], dotarray[119][4], dotarray[120][4], dotarray[121][4], dotarray[122][4], dotarray[123][4], dotarray[124][4], dotarray[125][4], dotarray[126][4], dotarray[127][4]};
assign dot_col_5 = {dotarray[0][5], dotarray[1][5], dotarray[2][5], dotarray[3][5], dotarray[4][5], dotarray[5][5], dotarray[6][5], dotarray[7][5], dotarray[8][5], dotarray[9][5], dotarray[10][5], dotarray[11][5], dotarray[12][5], dotarray[13][5], dotarray[14][5], dotarray[15][5], dotarray[16][5], dotarray[17][5], dotarray[18][5], dotarray[19][5], dotarray[20][5], dotarray[21][5], dotarray[22][5], dotarray[23][5], dotarray[24][5], dotarray[25][5], dotarray[26][5], dotarray[27][5], dotarray[28][5], dotarray[29][5], dotarray[30][5], dotarray[31][5], dotarray[32][5], dotarray[33][5], dotarray[34][5], dotarray[35][5], dotarray[36][5], dotarray[37][5], dotarray[38][5], dotarray[39][5], dotarray[40][5], dotarray[41][5], dotarray[42][5], dotarray[43][5], dotarray[44][5], dotarray[45][5], dotarray[46][5], dotarray[47][5], dotarray[48][5], dotarray[49][5], dotarray[50][5], dotarray[51][5], dotarray[52][5], dotarray[53][5], dotarray[54][5], dotarray[55][5], dotarray[56][5], dotarray[57][5], dotarray[58][5], dotarray[59][5], dotarray[60][5], dotarray[61][5], dotarray[62][5], dotarray[63][5], dotarray[64][5], dotarray[65][5], dotarray[66][5], dotarray[67][5], dotarray[68][5], dotarray[69][5], dotarray[70][5], dotarray[71][5], dotarray[72][5], dotarray[73][5], dotarray[74][5], dotarray[75][5], dotarray[76][5], dotarray[77][5], dotarray[78][5], dotarray[79][5], dotarray[80][5], dotarray[81][5], dotarray[82][5], dotarray[83][5], dotarray[84][5], dotarray[85][5], dotarray[86][5], dotarray[87][5], dotarray[88][5], dotarray[89][5], dotarray[90][5], dotarray[91][5], dotarray[92][5], dotarray[93][5], dotarray[94][5], dotarray[95][5], dotarray[96][5], dotarray[97][5], dotarray[98][5], dotarray[99][5], dotarray[100][5], dotarray[101][5], dotarray[102][5], dotarray[103][5], dotarray[104][5], dotarray[105][5], dotarray[106][5], dotarray[107][5], dotarray[108][5], dotarray[109][5], dotarray[110][5], dotarray[111][5], dotarray[112][5], dotarray[113][5], dotarray[114][5], dotarray[115][5], dotarray[116][5], dotarray[117][5], dotarray[118][5], dotarray[119][5], dotarray[120][5], dotarray[121][5], dotarray[122][5], dotarray[123][5], dotarray[124][5], dotarray[125][5], dotarray[126][5], dotarray[127][5]};
assign dot_col_6 = {dotarray[0][6], dotarray[1][6], dotarray[2][6], dotarray[3][6], dotarray[4][6], dotarray[5][6], dotarray[6][6], dotarray[7][6], dotarray[8][6], dotarray[9][6], dotarray[10][6], dotarray[11][6], dotarray[12][6], dotarray[13][6], dotarray[14][6], dotarray[15][6], dotarray[16][6], dotarray[17][6], dotarray[18][6], dotarray[19][6], dotarray[20][6], dotarray[21][6], dotarray[22][6], dotarray[23][6], dotarray[24][6], dotarray[25][6], dotarray[26][6], dotarray[27][6], dotarray[28][6], dotarray[29][6], dotarray[30][6], dotarray[31][6], dotarray[32][6], dotarray[33][6], dotarray[34][6], dotarray[35][6], dotarray[36][6], dotarray[37][6], dotarray[38][6], dotarray[39][6], dotarray[40][6], dotarray[41][6], dotarray[42][6], dotarray[43][6], dotarray[44][6], dotarray[45][6], dotarray[46][6], dotarray[47][6], dotarray[48][6], dotarray[49][6], dotarray[50][6], dotarray[51][6], dotarray[52][6], dotarray[53][6], dotarray[54][6], dotarray[55][6], dotarray[56][6], dotarray[57][6], dotarray[58][6], dotarray[59][6], dotarray[60][6], dotarray[61][6], dotarray[62][6], dotarray[63][6], dotarray[64][6], dotarray[65][6], dotarray[66][6], dotarray[67][6], dotarray[68][6], dotarray[69][6], dotarray[70][6], dotarray[71][6], dotarray[72][6], dotarray[73][6], dotarray[74][6], dotarray[75][6], dotarray[76][6], dotarray[77][6], dotarray[78][6], dotarray[79][6], dotarray[80][6], dotarray[81][6], dotarray[82][6], dotarray[83][6], dotarray[84][6], dotarray[85][6], dotarray[86][6], dotarray[87][6], dotarray[88][6], dotarray[89][6], dotarray[90][6], dotarray[91][6], dotarray[92][6], dotarray[93][6], dotarray[94][6], dotarray[95][6], dotarray[96][6], dotarray[97][6], dotarray[98][6], dotarray[99][6], dotarray[100][6], dotarray[101][6], dotarray[102][6], dotarray[103][6], dotarray[104][6], dotarray[105][6], dotarray[106][6], dotarray[107][6], dotarray[108][6], dotarray[109][6], dotarray[110][6], dotarray[111][6], dotarray[112][6], dotarray[113][6], dotarray[114][6], dotarray[115][6], dotarray[116][6], dotarray[117][6], dotarray[118][6], dotarray[119][6], dotarray[120][6], dotarray[121][6], dotarray[122][6], dotarray[123][6], dotarray[124][6], dotarray[125][6], dotarray[126][6], dotarray[127][6]};
assign dot_col_7 = {dotarray[0][7], dotarray[1][7], dotarray[2][7], dotarray[3][7], dotarray[4][7], dotarray[5][7], dotarray[6][7], dotarray[7][7], dotarray[8][7], dotarray[9][7], dotarray[10][7], dotarray[11][7], dotarray[12][7], dotarray[13][7], dotarray[14][7], dotarray[15][7], dotarray[16][7], dotarray[17][7], dotarray[18][7], dotarray[19][7], dotarray[20][7], dotarray[21][7], dotarray[22][7], dotarray[23][7], dotarray[24][7], dotarray[25][7], dotarray[26][7], dotarray[27][7], dotarray[28][7], dotarray[29][7], dotarray[30][7], dotarray[31][7], dotarray[32][7], dotarray[33][7], dotarray[34][7], dotarray[35][7], dotarray[36][7], dotarray[37][7], dotarray[38][7], dotarray[39][7], dotarray[40][7], dotarray[41][7], dotarray[42][7], dotarray[43][7], dotarray[44][7], dotarray[45][7], dotarray[46][7], dotarray[47][7], dotarray[48][7], dotarray[49][7], dotarray[50][7], dotarray[51][7], dotarray[52][7], dotarray[53][7], dotarray[54][7], dotarray[55][7], dotarray[56][7], dotarray[57][7], dotarray[58][7], dotarray[59][7], dotarray[60][7], dotarray[61][7], dotarray[62][7], dotarray[63][7], dotarray[64][7], dotarray[65][7], dotarray[66][7], dotarray[67][7], dotarray[68][7], dotarray[69][7], dotarray[70][7], dotarray[71][7], dotarray[72][7], dotarray[73][7], dotarray[74][7], dotarray[75][7], dotarray[76][7], dotarray[77][7], dotarray[78][7], dotarray[79][7], dotarray[80][7], dotarray[81][7], dotarray[82][7], dotarray[83][7], dotarray[84][7], dotarray[85][7], dotarray[86][7], dotarray[87][7], dotarray[88][7], dotarray[89][7], dotarray[90][7], dotarray[91][7], dotarray[92][7], dotarray[93][7], dotarray[94][7], dotarray[95][7], dotarray[96][7], dotarray[97][7], dotarray[98][7], dotarray[99][7], dotarray[100][7], dotarray[101][7], dotarray[102][7], dotarray[103][7], dotarray[104][7], dotarray[105][7], dotarray[106][7], dotarray[107][7], dotarray[108][7], dotarray[109][7], dotarray[110][7], dotarray[111][7], dotarray[112][7], dotarray[113][7], dotarray[114][7], dotarray[115][7], dotarray[116][7], dotarray[117][7], dotarray[118][7], dotarray[119][7], dotarray[120][7], dotarray[121][7], dotarray[122][7], dotarray[123][7], dotarray[124][7], dotarray[125][7], dotarray[126][7], dotarray[127][7]};
assign dot_col_8 = {dotarray[0][8], dotarray[1][8], dotarray[2][8], dotarray[3][8], dotarray[4][8], dotarray[5][8], dotarray[6][8], dotarray[7][8], dotarray[8][8], dotarray[9][8], dotarray[10][8], dotarray[11][8], dotarray[12][8], dotarray[13][8], dotarray[14][8], dotarray[15][8], dotarray[16][8], dotarray[17][8], dotarray[18][8], dotarray[19][8], dotarray[20][8], dotarray[21][8], dotarray[22][8], dotarray[23][8], dotarray[24][8], dotarray[25][8], dotarray[26][8], dotarray[27][8], dotarray[28][8], dotarray[29][8], dotarray[30][8], dotarray[31][8], dotarray[32][8], dotarray[33][8], dotarray[34][8], dotarray[35][8], dotarray[36][8], dotarray[37][8], dotarray[38][8], dotarray[39][8], dotarray[40][8], dotarray[41][8], dotarray[42][8], dotarray[43][8], dotarray[44][8], dotarray[45][8], dotarray[46][8], dotarray[47][8], dotarray[48][8], dotarray[49][8], dotarray[50][8], dotarray[51][8], dotarray[52][8], dotarray[53][8], dotarray[54][8], dotarray[55][8], dotarray[56][8], dotarray[57][8], dotarray[58][8], dotarray[59][8], dotarray[60][8], dotarray[61][8], dotarray[62][8], dotarray[63][8], dotarray[64][8], dotarray[65][8], dotarray[66][8], dotarray[67][8], dotarray[68][8], dotarray[69][8], dotarray[70][8], dotarray[71][8], dotarray[72][8], dotarray[73][8], dotarray[74][8], dotarray[75][8], dotarray[76][8], dotarray[77][8], dotarray[78][8], dotarray[79][8], dotarray[80][8], dotarray[81][8], dotarray[82][8], dotarray[83][8], dotarray[84][8], dotarray[85][8], dotarray[86][8], dotarray[87][8], dotarray[88][8], dotarray[89][8], dotarray[90][8], dotarray[91][8], dotarray[92][8], dotarray[93][8], dotarray[94][8], dotarray[95][8], dotarray[96][8], dotarray[97][8], dotarray[98][8], dotarray[99][8], dotarray[100][8], dotarray[101][8], dotarray[102][8], dotarray[103][8], dotarray[104][8], dotarray[105][8], dotarray[106][8], dotarray[107][8], dotarray[108][8], dotarray[109][8], dotarray[110][8], dotarray[111][8], dotarray[112][8], dotarray[113][8], dotarray[114][8], dotarray[115][8], dotarray[116][8], dotarray[117][8], dotarray[118][8], dotarray[119][8], dotarray[120][8], dotarray[121][8], dotarray[122][8], dotarray[123][8], dotarray[124][8], dotarray[125][8], dotarray[126][8], dotarray[127][8]};
assign dot_col_9 = {dotarray[0][9], dotarray[1][9], dotarray[2][9], dotarray[3][9], dotarray[4][9], dotarray[5][9], dotarray[6][9], dotarray[7][9], dotarray[8][9], dotarray[9][9], dotarray[10][9], dotarray[11][9], dotarray[12][9], dotarray[13][9], dotarray[14][9], dotarray[15][9], dotarray[16][9], dotarray[17][9], dotarray[18][9], dotarray[19][9], dotarray[20][9], dotarray[21][9], dotarray[22][9], dotarray[23][9], dotarray[24][9], dotarray[25][9], dotarray[26][9], dotarray[27][9], dotarray[28][9], dotarray[29][9], dotarray[30][9], dotarray[31][9], dotarray[32][9], dotarray[33][9], dotarray[34][9], dotarray[35][9], dotarray[36][9], dotarray[37][9], dotarray[38][9], dotarray[39][9], dotarray[40][9], dotarray[41][9], dotarray[42][9], dotarray[43][9], dotarray[44][9], dotarray[45][9], dotarray[46][9], dotarray[47][9], dotarray[48][9], dotarray[49][9], dotarray[50][9], dotarray[51][9], dotarray[52][9], dotarray[53][9], dotarray[54][9], dotarray[55][9], dotarray[56][9], dotarray[57][9], dotarray[58][9], dotarray[59][9], dotarray[60][9], dotarray[61][9], dotarray[62][9], dotarray[63][9], dotarray[64][9], dotarray[65][9], dotarray[66][9], dotarray[67][9], dotarray[68][9], dotarray[69][9], dotarray[70][9], dotarray[71][9], dotarray[72][9], dotarray[73][9], dotarray[74][9], dotarray[75][9], dotarray[76][9], dotarray[77][9], dotarray[78][9], dotarray[79][9], dotarray[80][9], dotarray[81][9], dotarray[82][9], dotarray[83][9], dotarray[84][9], dotarray[85][9], dotarray[86][9], dotarray[87][9], dotarray[88][9], dotarray[89][9], dotarray[90][9], dotarray[91][9], dotarray[92][9], dotarray[93][9], dotarray[94][9], dotarray[95][9], dotarray[96][9], dotarray[97][9], dotarray[98][9], dotarray[99][9], dotarray[100][9], dotarray[101][9], dotarray[102][9], dotarray[103][9], dotarray[104][9], dotarray[105][9], dotarray[106][9], dotarray[107][9], dotarray[108][9], dotarray[109][9], dotarray[110][9], dotarray[111][9], dotarray[112][9], dotarray[113][9], dotarray[114][9], dotarray[115][9], dotarray[116][9], dotarray[117][9], dotarray[118][9], dotarray[119][9], dotarray[120][9], dotarray[121][9], dotarray[122][9], dotarray[123][9], dotarray[124][9], dotarray[125][9], dotarray[126][9], dotarray[127][9]};
assign dot_col_10 = {dotarray[0][10], dotarray[1][10], dotarray[2][10], dotarray[3][10], dotarray[4][10], dotarray[5][10], dotarray[6][10], dotarray[7][10], dotarray[8][10], dotarray[9][10], dotarray[10][10], dotarray[11][10], dotarray[12][10], dotarray[13][10], dotarray[14][10], dotarray[15][10], dotarray[16][10], dotarray[17][10], dotarray[18][10], dotarray[19][10], dotarray[20][10], dotarray[21][10], dotarray[22][10], dotarray[23][10], dotarray[24][10], dotarray[25][10], dotarray[26][10], dotarray[27][10], dotarray[28][10], dotarray[29][10], dotarray[30][10], dotarray[31][10], dotarray[32][10], dotarray[33][10], dotarray[34][10], dotarray[35][10], dotarray[36][10], dotarray[37][10], dotarray[38][10], dotarray[39][10], dotarray[40][10], dotarray[41][10], dotarray[42][10], dotarray[43][10], dotarray[44][10], dotarray[45][10], dotarray[46][10], dotarray[47][10], dotarray[48][10], dotarray[49][10], dotarray[50][10], dotarray[51][10], dotarray[52][10], dotarray[53][10], dotarray[54][10], dotarray[55][10], dotarray[56][10], dotarray[57][10], dotarray[58][10], dotarray[59][10], dotarray[60][10], dotarray[61][10], dotarray[62][10], dotarray[63][10], dotarray[64][10], dotarray[65][10], dotarray[66][10], dotarray[67][10], dotarray[68][10], dotarray[69][10], dotarray[70][10], dotarray[71][10], dotarray[72][10], dotarray[73][10], dotarray[74][10], dotarray[75][10], dotarray[76][10], dotarray[77][10], dotarray[78][10], dotarray[79][10], dotarray[80][10], dotarray[81][10], dotarray[82][10], dotarray[83][10], dotarray[84][10], dotarray[85][10], dotarray[86][10], dotarray[87][10], dotarray[88][10], dotarray[89][10], dotarray[90][10], dotarray[91][10], dotarray[92][10], dotarray[93][10], dotarray[94][10], dotarray[95][10], dotarray[96][10], dotarray[97][10], dotarray[98][10], dotarray[99][10], dotarray[100][10], dotarray[101][10], dotarray[102][10], dotarray[103][10], dotarray[104][10], dotarray[105][10], dotarray[106][10], dotarray[107][10], dotarray[108][10], dotarray[109][10], dotarray[110][10], dotarray[111][10], dotarray[112][10], dotarray[113][10], dotarray[114][10], dotarray[115][10], dotarray[116][10], dotarray[117][10], dotarray[118][10], dotarray[119][10], dotarray[120][10], dotarray[121][10], dotarray[122][10], dotarray[123][10], dotarray[124][10], dotarray[125][10], dotarray[126][10], dotarray[127][10]};
assign dot_col_11 = {dotarray[0][11], dotarray[1][11], dotarray[2][11], dotarray[3][11], dotarray[4][11], dotarray[5][11], dotarray[6][11], dotarray[7][11], dotarray[8][11], dotarray[9][11], dotarray[10][11], dotarray[11][11], dotarray[12][11], dotarray[13][11], dotarray[14][11], dotarray[15][11], dotarray[16][11], dotarray[17][11], dotarray[18][11], dotarray[19][11], dotarray[20][11], dotarray[21][11], dotarray[22][11], dotarray[23][11], dotarray[24][11], dotarray[25][11], dotarray[26][11], dotarray[27][11], dotarray[28][11], dotarray[29][11], dotarray[30][11], dotarray[31][11], dotarray[32][11], dotarray[33][11], dotarray[34][11], dotarray[35][11], dotarray[36][11], dotarray[37][11], dotarray[38][11], dotarray[39][11], dotarray[40][11], dotarray[41][11], dotarray[42][11], dotarray[43][11], dotarray[44][11], dotarray[45][11], dotarray[46][11], dotarray[47][11], dotarray[48][11], dotarray[49][11], dotarray[50][11], dotarray[51][11], dotarray[52][11], dotarray[53][11], dotarray[54][11], dotarray[55][11], dotarray[56][11], dotarray[57][11], dotarray[58][11], dotarray[59][11], dotarray[60][11], dotarray[61][11], dotarray[62][11], dotarray[63][11], dotarray[64][11], dotarray[65][11], dotarray[66][11], dotarray[67][11], dotarray[68][11], dotarray[69][11], dotarray[70][11], dotarray[71][11], dotarray[72][11], dotarray[73][11], dotarray[74][11], dotarray[75][11], dotarray[76][11], dotarray[77][11], dotarray[78][11], dotarray[79][11], dotarray[80][11], dotarray[81][11], dotarray[82][11], dotarray[83][11], dotarray[84][11], dotarray[85][11], dotarray[86][11], dotarray[87][11], dotarray[88][11], dotarray[89][11], dotarray[90][11], dotarray[91][11], dotarray[92][11], dotarray[93][11], dotarray[94][11], dotarray[95][11], dotarray[96][11], dotarray[97][11], dotarray[98][11], dotarray[99][11], dotarray[100][11], dotarray[101][11], dotarray[102][11], dotarray[103][11], dotarray[104][11], dotarray[105][11], dotarray[106][11], dotarray[107][11], dotarray[108][11], dotarray[109][11], dotarray[110][11], dotarray[111][11], dotarray[112][11], dotarray[113][11], dotarray[114][11], dotarray[115][11], dotarray[116][11], dotarray[117][11], dotarray[118][11], dotarray[119][11], dotarray[120][11], dotarray[121][11], dotarray[122][11], dotarray[123][11], dotarray[124][11], dotarray[125][11], dotarray[126][11], dotarray[127][11]};
assign dot_col_12 = {dotarray[0][12], dotarray[1][12], dotarray[2][12], dotarray[3][12], dotarray[4][12], dotarray[5][12], dotarray[6][12], dotarray[7][12], dotarray[8][12], dotarray[9][12], dotarray[10][12], dotarray[11][12], dotarray[12][12], dotarray[13][12], dotarray[14][12], dotarray[15][12], dotarray[16][12], dotarray[17][12], dotarray[18][12], dotarray[19][12], dotarray[20][12], dotarray[21][12], dotarray[22][12], dotarray[23][12], dotarray[24][12], dotarray[25][12], dotarray[26][12], dotarray[27][12], dotarray[28][12], dotarray[29][12], dotarray[30][12], dotarray[31][12], dotarray[32][12], dotarray[33][12], dotarray[34][12], dotarray[35][12], dotarray[36][12], dotarray[37][12], dotarray[38][12], dotarray[39][12], dotarray[40][12], dotarray[41][12], dotarray[42][12], dotarray[43][12], dotarray[44][12], dotarray[45][12], dotarray[46][12], dotarray[47][12], dotarray[48][12], dotarray[49][12], dotarray[50][12], dotarray[51][12], dotarray[52][12], dotarray[53][12], dotarray[54][12], dotarray[55][12], dotarray[56][12], dotarray[57][12], dotarray[58][12], dotarray[59][12], dotarray[60][12], dotarray[61][12], dotarray[62][12], dotarray[63][12], dotarray[64][12], dotarray[65][12], dotarray[66][12], dotarray[67][12], dotarray[68][12], dotarray[69][12], dotarray[70][12], dotarray[71][12], dotarray[72][12], dotarray[73][12], dotarray[74][12], dotarray[75][12], dotarray[76][12], dotarray[77][12], dotarray[78][12], dotarray[79][12], dotarray[80][12], dotarray[81][12], dotarray[82][12], dotarray[83][12], dotarray[84][12], dotarray[85][12], dotarray[86][12], dotarray[87][12], dotarray[88][12], dotarray[89][12], dotarray[90][12], dotarray[91][12], dotarray[92][12], dotarray[93][12], dotarray[94][12], dotarray[95][12], dotarray[96][12], dotarray[97][12], dotarray[98][12], dotarray[99][12], dotarray[100][12], dotarray[101][12], dotarray[102][12], dotarray[103][12], dotarray[104][12], dotarray[105][12], dotarray[106][12], dotarray[107][12], dotarray[108][12], dotarray[109][12], dotarray[110][12], dotarray[111][12], dotarray[112][12], dotarray[113][12], dotarray[114][12], dotarray[115][12], dotarray[116][12], dotarray[117][12], dotarray[118][12], dotarray[119][12], dotarray[120][12], dotarray[121][12], dotarray[122][12], dotarray[123][12], dotarray[124][12], dotarray[125][12], dotarray[126][12], dotarray[127][12]};
assign dot_col_13 = {dotarray[0][13], dotarray[1][13], dotarray[2][13], dotarray[3][13], dotarray[4][13], dotarray[5][13], dotarray[6][13], dotarray[7][13], dotarray[8][13], dotarray[9][13], dotarray[10][13], dotarray[11][13], dotarray[12][13], dotarray[13][13], dotarray[14][13], dotarray[15][13], dotarray[16][13], dotarray[17][13], dotarray[18][13], dotarray[19][13], dotarray[20][13], dotarray[21][13], dotarray[22][13], dotarray[23][13], dotarray[24][13], dotarray[25][13], dotarray[26][13], dotarray[27][13], dotarray[28][13], dotarray[29][13], dotarray[30][13], dotarray[31][13], dotarray[32][13], dotarray[33][13], dotarray[34][13], dotarray[35][13], dotarray[36][13], dotarray[37][13], dotarray[38][13], dotarray[39][13], dotarray[40][13], dotarray[41][13], dotarray[42][13], dotarray[43][13], dotarray[44][13], dotarray[45][13], dotarray[46][13], dotarray[47][13], dotarray[48][13], dotarray[49][13], dotarray[50][13], dotarray[51][13], dotarray[52][13], dotarray[53][13], dotarray[54][13], dotarray[55][13], dotarray[56][13], dotarray[57][13], dotarray[58][13], dotarray[59][13], dotarray[60][13], dotarray[61][13], dotarray[62][13], dotarray[63][13], dotarray[64][13], dotarray[65][13], dotarray[66][13], dotarray[67][13], dotarray[68][13], dotarray[69][13], dotarray[70][13], dotarray[71][13], dotarray[72][13], dotarray[73][13], dotarray[74][13], dotarray[75][13], dotarray[76][13], dotarray[77][13], dotarray[78][13], dotarray[79][13], dotarray[80][13], dotarray[81][13], dotarray[82][13], dotarray[83][13], dotarray[84][13], dotarray[85][13], dotarray[86][13], dotarray[87][13], dotarray[88][13], dotarray[89][13], dotarray[90][13], dotarray[91][13], dotarray[92][13], dotarray[93][13], dotarray[94][13], dotarray[95][13], dotarray[96][13], dotarray[97][13], dotarray[98][13], dotarray[99][13], dotarray[100][13], dotarray[101][13], dotarray[102][13], dotarray[103][13], dotarray[104][13], dotarray[105][13], dotarray[106][13], dotarray[107][13], dotarray[108][13], dotarray[109][13], dotarray[110][13], dotarray[111][13], dotarray[112][13], dotarray[113][13], dotarray[114][13], dotarray[115][13], dotarray[116][13], dotarray[117][13], dotarray[118][13], dotarray[119][13], dotarray[120][13], dotarray[121][13], dotarray[122][13], dotarray[123][13], dotarray[124][13], dotarray[125][13], dotarray[126][13], dotarray[127][13]};
assign dot_col_14 = {dotarray[0][14], dotarray[1][14], dotarray[2][14], dotarray[3][14], dotarray[4][14], dotarray[5][14], dotarray[6][14], dotarray[7][14], dotarray[8][14], dotarray[9][14], dotarray[10][14], dotarray[11][14], dotarray[12][14], dotarray[13][14], dotarray[14][14], dotarray[15][14], dotarray[16][14], dotarray[17][14], dotarray[18][14], dotarray[19][14], dotarray[20][14], dotarray[21][14], dotarray[22][14], dotarray[23][14], dotarray[24][14], dotarray[25][14], dotarray[26][14], dotarray[27][14], dotarray[28][14], dotarray[29][14], dotarray[30][14], dotarray[31][14], dotarray[32][14], dotarray[33][14], dotarray[34][14], dotarray[35][14], dotarray[36][14], dotarray[37][14], dotarray[38][14], dotarray[39][14], dotarray[40][14], dotarray[41][14], dotarray[42][14], dotarray[43][14], dotarray[44][14], dotarray[45][14], dotarray[46][14], dotarray[47][14], dotarray[48][14], dotarray[49][14], dotarray[50][14], dotarray[51][14], dotarray[52][14], dotarray[53][14], dotarray[54][14], dotarray[55][14], dotarray[56][14], dotarray[57][14], dotarray[58][14], dotarray[59][14], dotarray[60][14], dotarray[61][14], dotarray[62][14], dotarray[63][14], dotarray[64][14], dotarray[65][14], dotarray[66][14], dotarray[67][14], dotarray[68][14], dotarray[69][14], dotarray[70][14], dotarray[71][14], dotarray[72][14], dotarray[73][14], dotarray[74][14], dotarray[75][14], dotarray[76][14], dotarray[77][14], dotarray[78][14], dotarray[79][14], dotarray[80][14], dotarray[81][14], dotarray[82][14], dotarray[83][14], dotarray[84][14], dotarray[85][14], dotarray[86][14], dotarray[87][14], dotarray[88][14], dotarray[89][14], dotarray[90][14], dotarray[91][14], dotarray[92][14], dotarray[93][14], dotarray[94][14], dotarray[95][14], dotarray[96][14], dotarray[97][14], dotarray[98][14], dotarray[99][14], dotarray[100][14], dotarray[101][14], dotarray[102][14], dotarray[103][14], dotarray[104][14], dotarray[105][14], dotarray[106][14], dotarray[107][14], dotarray[108][14], dotarray[109][14], dotarray[110][14], dotarray[111][14], dotarray[112][14], dotarray[113][14], dotarray[114][14], dotarray[115][14], dotarray[116][14], dotarray[117][14], dotarray[118][14], dotarray[119][14], dotarray[120][14], dotarray[121][14], dotarray[122][14], dotarray[123][14], dotarray[124][14], dotarray[125][14], dotarray[126][14], dotarray[127][14]};
assign dot_col_15 = {dotarray[0][15], dotarray[1][15], dotarray[2][15], dotarray[3][15], dotarray[4][15], dotarray[5][15], dotarray[6][15], dotarray[7][15], dotarray[8][15], dotarray[9][15], dotarray[10][15], dotarray[11][15], dotarray[12][15], dotarray[13][15], dotarray[14][15], dotarray[15][15], dotarray[16][15], dotarray[17][15], dotarray[18][15], dotarray[19][15], dotarray[20][15], dotarray[21][15], dotarray[22][15], dotarray[23][15], dotarray[24][15], dotarray[25][15], dotarray[26][15], dotarray[27][15], dotarray[28][15], dotarray[29][15], dotarray[30][15], dotarray[31][15], dotarray[32][15], dotarray[33][15], dotarray[34][15], dotarray[35][15], dotarray[36][15], dotarray[37][15], dotarray[38][15], dotarray[39][15], dotarray[40][15], dotarray[41][15], dotarray[42][15], dotarray[43][15], dotarray[44][15], dotarray[45][15], dotarray[46][15], dotarray[47][15], dotarray[48][15], dotarray[49][15], dotarray[50][15], dotarray[51][15], dotarray[52][15], dotarray[53][15], dotarray[54][15], dotarray[55][15], dotarray[56][15], dotarray[57][15], dotarray[58][15], dotarray[59][15], dotarray[60][15], dotarray[61][15], dotarray[62][15], dotarray[63][15], dotarray[64][15], dotarray[65][15], dotarray[66][15], dotarray[67][15], dotarray[68][15], dotarray[69][15], dotarray[70][15], dotarray[71][15], dotarray[72][15], dotarray[73][15], dotarray[74][15], dotarray[75][15], dotarray[76][15], dotarray[77][15], dotarray[78][15], dotarray[79][15], dotarray[80][15], dotarray[81][15], dotarray[82][15], dotarray[83][15], dotarray[84][15], dotarray[85][15], dotarray[86][15], dotarray[87][15], dotarray[88][15], dotarray[89][15], dotarray[90][15], dotarray[91][15], dotarray[92][15], dotarray[93][15], dotarray[94][15], dotarray[95][15], dotarray[96][15], dotarray[97][15], dotarray[98][15], dotarray[99][15], dotarray[100][15], dotarray[101][15], dotarray[102][15], dotarray[103][15], dotarray[104][15], dotarray[105][15], dotarray[106][15], dotarray[107][15], dotarray[108][15], dotarray[109][15], dotarray[110][15], dotarray[111][15], dotarray[112][15], dotarray[113][15], dotarray[114][15], dotarray[115][15], dotarray[116][15], dotarray[117][15], dotarray[118][15], dotarray[119][15], dotarray[120][15], dotarray[121][15], dotarray[122][15], dotarray[123][15], dotarray[124][15], dotarray[125][15], dotarray[126][15], dotarray[127][15]};
assign dot_col_16 = {dotarray[0][16], dotarray[1][16], dotarray[2][16], dotarray[3][16], dotarray[4][16], dotarray[5][16], dotarray[6][16], dotarray[7][16], dotarray[8][16], dotarray[9][16], dotarray[10][16], dotarray[11][16], dotarray[12][16], dotarray[13][16], dotarray[14][16], dotarray[15][16], dotarray[16][16], dotarray[17][16], dotarray[18][16], dotarray[19][16], dotarray[20][16], dotarray[21][16], dotarray[22][16], dotarray[23][16], dotarray[24][16], dotarray[25][16], dotarray[26][16], dotarray[27][16], dotarray[28][16], dotarray[29][16], dotarray[30][16], dotarray[31][16], dotarray[32][16], dotarray[33][16], dotarray[34][16], dotarray[35][16], dotarray[36][16], dotarray[37][16], dotarray[38][16], dotarray[39][16], dotarray[40][16], dotarray[41][16], dotarray[42][16], dotarray[43][16], dotarray[44][16], dotarray[45][16], dotarray[46][16], dotarray[47][16], dotarray[48][16], dotarray[49][16], dotarray[50][16], dotarray[51][16], dotarray[52][16], dotarray[53][16], dotarray[54][16], dotarray[55][16], dotarray[56][16], dotarray[57][16], dotarray[58][16], dotarray[59][16], dotarray[60][16], dotarray[61][16], dotarray[62][16], dotarray[63][16], dotarray[64][16], dotarray[65][16], dotarray[66][16], dotarray[67][16], dotarray[68][16], dotarray[69][16], dotarray[70][16], dotarray[71][16], dotarray[72][16], dotarray[73][16], dotarray[74][16], dotarray[75][16], dotarray[76][16], dotarray[77][16], dotarray[78][16], dotarray[79][16], dotarray[80][16], dotarray[81][16], dotarray[82][16], dotarray[83][16], dotarray[84][16], dotarray[85][16], dotarray[86][16], dotarray[87][16], dotarray[88][16], dotarray[89][16], dotarray[90][16], dotarray[91][16], dotarray[92][16], dotarray[93][16], dotarray[94][16], dotarray[95][16], dotarray[96][16], dotarray[97][16], dotarray[98][16], dotarray[99][16], dotarray[100][16], dotarray[101][16], dotarray[102][16], dotarray[103][16], dotarray[104][16], dotarray[105][16], dotarray[106][16], dotarray[107][16], dotarray[108][16], dotarray[109][16], dotarray[110][16], dotarray[111][16], dotarray[112][16], dotarray[113][16], dotarray[114][16], dotarray[115][16], dotarray[116][16], dotarray[117][16], dotarray[118][16], dotarray[119][16], dotarray[120][16], dotarray[121][16], dotarray[122][16], dotarray[123][16], dotarray[124][16], dotarray[125][16], dotarray[126][16], dotarray[127][16]};
assign dot_col_17 = {dotarray[0][17], dotarray[1][17], dotarray[2][17], dotarray[3][17], dotarray[4][17], dotarray[5][17], dotarray[6][17], dotarray[7][17], dotarray[8][17], dotarray[9][17], dotarray[10][17], dotarray[11][17], dotarray[12][17], dotarray[13][17], dotarray[14][17], dotarray[15][17], dotarray[16][17], dotarray[17][17], dotarray[18][17], dotarray[19][17], dotarray[20][17], dotarray[21][17], dotarray[22][17], dotarray[23][17], dotarray[24][17], dotarray[25][17], dotarray[26][17], dotarray[27][17], dotarray[28][17], dotarray[29][17], dotarray[30][17], dotarray[31][17], dotarray[32][17], dotarray[33][17], dotarray[34][17], dotarray[35][17], dotarray[36][17], dotarray[37][17], dotarray[38][17], dotarray[39][17], dotarray[40][17], dotarray[41][17], dotarray[42][17], dotarray[43][17], dotarray[44][17], dotarray[45][17], dotarray[46][17], dotarray[47][17], dotarray[48][17], dotarray[49][17], dotarray[50][17], dotarray[51][17], dotarray[52][17], dotarray[53][17], dotarray[54][17], dotarray[55][17], dotarray[56][17], dotarray[57][17], dotarray[58][17], dotarray[59][17], dotarray[60][17], dotarray[61][17], dotarray[62][17], dotarray[63][17], dotarray[64][17], dotarray[65][17], dotarray[66][17], dotarray[67][17], dotarray[68][17], dotarray[69][17], dotarray[70][17], dotarray[71][17], dotarray[72][17], dotarray[73][17], dotarray[74][17], dotarray[75][17], dotarray[76][17], dotarray[77][17], dotarray[78][17], dotarray[79][17], dotarray[80][17], dotarray[81][17], dotarray[82][17], dotarray[83][17], dotarray[84][17], dotarray[85][17], dotarray[86][17], dotarray[87][17], dotarray[88][17], dotarray[89][17], dotarray[90][17], dotarray[91][17], dotarray[92][17], dotarray[93][17], dotarray[94][17], dotarray[95][17], dotarray[96][17], dotarray[97][17], dotarray[98][17], dotarray[99][17], dotarray[100][17], dotarray[101][17], dotarray[102][17], dotarray[103][17], dotarray[104][17], dotarray[105][17], dotarray[106][17], dotarray[107][17], dotarray[108][17], dotarray[109][17], dotarray[110][17], dotarray[111][17], dotarray[112][17], dotarray[113][17], dotarray[114][17], dotarray[115][17], dotarray[116][17], dotarray[117][17], dotarray[118][17], dotarray[119][17], dotarray[120][17], dotarray[121][17], dotarray[122][17], dotarray[123][17], dotarray[124][17], dotarray[125][17], dotarray[126][17], dotarray[127][17]};
assign dot_col_18 = {dotarray[0][18], dotarray[1][18], dotarray[2][18], dotarray[3][18], dotarray[4][18], dotarray[5][18], dotarray[6][18], dotarray[7][18], dotarray[8][18], dotarray[9][18], dotarray[10][18], dotarray[11][18], dotarray[12][18], dotarray[13][18], dotarray[14][18], dotarray[15][18], dotarray[16][18], dotarray[17][18], dotarray[18][18], dotarray[19][18], dotarray[20][18], dotarray[21][18], dotarray[22][18], dotarray[23][18], dotarray[24][18], dotarray[25][18], dotarray[26][18], dotarray[27][18], dotarray[28][18], dotarray[29][18], dotarray[30][18], dotarray[31][18], dotarray[32][18], dotarray[33][18], dotarray[34][18], dotarray[35][18], dotarray[36][18], dotarray[37][18], dotarray[38][18], dotarray[39][18], dotarray[40][18], dotarray[41][18], dotarray[42][18], dotarray[43][18], dotarray[44][18], dotarray[45][18], dotarray[46][18], dotarray[47][18], dotarray[48][18], dotarray[49][18], dotarray[50][18], dotarray[51][18], dotarray[52][18], dotarray[53][18], dotarray[54][18], dotarray[55][18], dotarray[56][18], dotarray[57][18], dotarray[58][18], dotarray[59][18], dotarray[60][18], dotarray[61][18], dotarray[62][18], dotarray[63][18], dotarray[64][18], dotarray[65][18], dotarray[66][18], dotarray[67][18], dotarray[68][18], dotarray[69][18], dotarray[70][18], dotarray[71][18], dotarray[72][18], dotarray[73][18], dotarray[74][18], dotarray[75][18], dotarray[76][18], dotarray[77][18], dotarray[78][18], dotarray[79][18], dotarray[80][18], dotarray[81][18], dotarray[82][18], dotarray[83][18], dotarray[84][18], dotarray[85][18], dotarray[86][18], dotarray[87][18], dotarray[88][18], dotarray[89][18], dotarray[90][18], dotarray[91][18], dotarray[92][18], dotarray[93][18], dotarray[94][18], dotarray[95][18], dotarray[96][18], dotarray[97][18], dotarray[98][18], dotarray[99][18], dotarray[100][18], dotarray[101][18], dotarray[102][18], dotarray[103][18], dotarray[104][18], dotarray[105][18], dotarray[106][18], dotarray[107][18], dotarray[108][18], dotarray[109][18], dotarray[110][18], dotarray[111][18], dotarray[112][18], dotarray[113][18], dotarray[114][18], dotarray[115][18], dotarray[116][18], dotarray[117][18], dotarray[118][18], dotarray[119][18], dotarray[120][18], dotarray[121][18], dotarray[122][18], dotarray[123][18], dotarray[124][18], dotarray[125][18], dotarray[126][18], dotarray[127][18]};
assign dot_col_19 = {dotarray[0][19], dotarray[1][19], dotarray[2][19], dotarray[3][19], dotarray[4][19], dotarray[5][19], dotarray[6][19], dotarray[7][19], dotarray[8][19], dotarray[9][19], dotarray[10][19], dotarray[11][19], dotarray[12][19], dotarray[13][19], dotarray[14][19], dotarray[15][19], dotarray[16][19], dotarray[17][19], dotarray[18][19], dotarray[19][19], dotarray[20][19], dotarray[21][19], dotarray[22][19], dotarray[23][19], dotarray[24][19], dotarray[25][19], dotarray[26][19], dotarray[27][19], dotarray[28][19], dotarray[29][19], dotarray[30][19], dotarray[31][19], dotarray[32][19], dotarray[33][19], dotarray[34][19], dotarray[35][19], dotarray[36][19], dotarray[37][19], dotarray[38][19], dotarray[39][19], dotarray[40][19], dotarray[41][19], dotarray[42][19], dotarray[43][19], dotarray[44][19], dotarray[45][19], dotarray[46][19], dotarray[47][19], dotarray[48][19], dotarray[49][19], dotarray[50][19], dotarray[51][19], dotarray[52][19], dotarray[53][19], dotarray[54][19], dotarray[55][19], dotarray[56][19], dotarray[57][19], dotarray[58][19], dotarray[59][19], dotarray[60][19], dotarray[61][19], dotarray[62][19], dotarray[63][19], dotarray[64][19], dotarray[65][19], dotarray[66][19], dotarray[67][19], dotarray[68][19], dotarray[69][19], dotarray[70][19], dotarray[71][19], dotarray[72][19], dotarray[73][19], dotarray[74][19], dotarray[75][19], dotarray[76][19], dotarray[77][19], dotarray[78][19], dotarray[79][19], dotarray[80][19], dotarray[81][19], dotarray[82][19], dotarray[83][19], dotarray[84][19], dotarray[85][19], dotarray[86][19], dotarray[87][19], dotarray[88][19], dotarray[89][19], dotarray[90][19], dotarray[91][19], dotarray[92][19], dotarray[93][19], dotarray[94][19], dotarray[95][19], dotarray[96][19], dotarray[97][19], dotarray[98][19], dotarray[99][19], dotarray[100][19], dotarray[101][19], dotarray[102][19], dotarray[103][19], dotarray[104][19], dotarray[105][19], dotarray[106][19], dotarray[107][19], dotarray[108][19], dotarray[109][19], dotarray[110][19], dotarray[111][19], dotarray[112][19], dotarray[113][19], dotarray[114][19], dotarray[115][19], dotarray[116][19], dotarray[117][19], dotarray[118][19], dotarray[119][19], dotarray[120][19], dotarray[121][19], dotarray[122][19], dotarray[123][19], dotarray[124][19], dotarray[125][19], dotarray[126][19], dotarray[127][19]};
assign dot_col_20 = {dotarray[0][20], dotarray[1][20], dotarray[2][20], dotarray[3][20], dotarray[4][20], dotarray[5][20], dotarray[6][20], dotarray[7][20], dotarray[8][20], dotarray[9][20], dotarray[10][20], dotarray[11][20], dotarray[12][20], dotarray[13][20], dotarray[14][20], dotarray[15][20], dotarray[16][20], dotarray[17][20], dotarray[18][20], dotarray[19][20], dotarray[20][20], dotarray[21][20], dotarray[22][20], dotarray[23][20], dotarray[24][20], dotarray[25][20], dotarray[26][20], dotarray[27][20], dotarray[28][20], dotarray[29][20], dotarray[30][20], dotarray[31][20], dotarray[32][20], dotarray[33][20], dotarray[34][20], dotarray[35][20], dotarray[36][20], dotarray[37][20], dotarray[38][20], dotarray[39][20], dotarray[40][20], dotarray[41][20], dotarray[42][20], dotarray[43][20], dotarray[44][20], dotarray[45][20], dotarray[46][20], dotarray[47][20], dotarray[48][20], dotarray[49][20], dotarray[50][20], dotarray[51][20], dotarray[52][20], dotarray[53][20], dotarray[54][20], dotarray[55][20], dotarray[56][20], dotarray[57][20], dotarray[58][20], dotarray[59][20], dotarray[60][20], dotarray[61][20], dotarray[62][20], dotarray[63][20], dotarray[64][20], dotarray[65][20], dotarray[66][20], dotarray[67][20], dotarray[68][20], dotarray[69][20], dotarray[70][20], dotarray[71][20], dotarray[72][20], dotarray[73][20], dotarray[74][20], dotarray[75][20], dotarray[76][20], dotarray[77][20], dotarray[78][20], dotarray[79][20], dotarray[80][20], dotarray[81][20], dotarray[82][20], dotarray[83][20], dotarray[84][20], dotarray[85][20], dotarray[86][20], dotarray[87][20], dotarray[88][20], dotarray[89][20], dotarray[90][20], dotarray[91][20], dotarray[92][20], dotarray[93][20], dotarray[94][20], dotarray[95][20], dotarray[96][20], dotarray[97][20], dotarray[98][20], dotarray[99][20], dotarray[100][20], dotarray[101][20], dotarray[102][20], dotarray[103][20], dotarray[104][20], dotarray[105][20], dotarray[106][20], dotarray[107][20], dotarray[108][20], dotarray[109][20], dotarray[110][20], dotarray[111][20], dotarray[112][20], dotarray[113][20], dotarray[114][20], dotarray[115][20], dotarray[116][20], dotarray[117][20], dotarray[118][20], dotarray[119][20], dotarray[120][20], dotarray[121][20], dotarray[122][20], dotarray[123][20], dotarray[124][20], dotarray[125][20], dotarray[126][20], dotarray[127][20]};
assign dot_col_21 = {dotarray[0][21], dotarray[1][21], dotarray[2][21], dotarray[3][21], dotarray[4][21], dotarray[5][21], dotarray[6][21], dotarray[7][21], dotarray[8][21], dotarray[9][21], dotarray[10][21], dotarray[11][21], dotarray[12][21], dotarray[13][21], dotarray[14][21], dotarray[15][21], dotarray[16][21], dotarray[17][21], dotarray[18][21], dotarray[19][21], dotarray[20][21], dotarray[21][21], dotarray[22][21], dotarray[23][21], dotarray[24][21], dotarray[25][21], dotarray[26][21], dotarray[27][21], dotarray[28][21], dotarray[29][21], dotarray[30][21], dotarray[31][21], dotarray[32][21], dotarray[33][21], dotarray[34][21], dotarray[35][21], dotarray[36][21], dotarray[37][21], dotarray[38][21], dotarray[39][21], dotarray[40][21], dotarray[41][21], dotarray[42][21], dotarray[43][21], dotarray[44][21], dotarray[45][21], dotarray[46][21], dotarray[47][21], dotarray[48][21], dotarray[49][21], dotarray[50][21], dotarray[51][21], dotarray[52][21], dotarray[53][21], dotarray[54][21], dotarray[55][21], dotarray[56][21], dotarray[57][21], dotarray[58][21], dotarray[59][21], dotarray[60][21], dotarray[61][21], dotarray[62][21], dotarray[63][21], dotarray[64][21], dotarray[65][21], dotarray[66][21], dotarray[67][21], dotarray[68][21], dotarray[69][21], dotarray[70][21], dotarray[71][21], dotarray[72][21], dotarray[73][21], dotarray[74][21], dotarray[75][21], dotarray[76][21], dotarray[77][21], dotarray[78][21], dotarray[79][21], dotarray[80][21], dotarray[81][21], dotarray[82][21], dotarray[83][21], dotarray[84][21], dotarray[85][21], dotarray[86][21], dotarray[87][21], dotarray[88][21], dotarray[89][21], dotarray[90][21], dotarray[91][21], dotarray[92][21], dotarray[93][21], dotarray[94][21], dotarray[95][21], dotarray[96][21], dotarray[97][21], dotarray[98][21], dotarray[99][21], dotarray[100][21], dotarray[101][21], dotarray[102][21], dotarray[103][21], dotarray[104][21], dotarray[105][21], dotarray[106][21], dotarray[107][21], dotarray[108][21], dotarray[109][21], dotarray[110][21], dotarray[111][21], dotarray[112][21], dotarray[113][21], dotarray[114][21], dotarray[115][21], dotarray[116][21], dotarray[117][21], dotarray[118][21], dotarray[119][21], dotarray[120][21], dotarray[121][21], dotarray[122][21], dotarray[123][21], dotarray[124][21], dotarray[125][21], dotarray[126][21], dotarray[127][21]};
assign dot_col_22 = {dotarray[0][22], dotarray[1][22], dotarray[2][22], dotarray[3][22], dotarray[4][22], dotarray[5][22], dotarray[6][22], dotarray[7][22], dotarray[8][22], dotarray[9][22], dotarray[10][22], dotarray[11][22], dotarray[12][22], dotarray[13][22], dotarray[14][22], dotarray[15][22], dotarray[16][22], dotarray[17][22], dotarray[18][22], dotarray[19][22], dotarray[20][22], dotarray[21][22], dotarray[22][22], dotarray[23][22], dotarray[24][22], dotarray[25][22], dotarray[26][22], dotarray[27][22], dotarray[28][22], dotarray[29][22], dotarray[30][22], dotarray[31][22], dotarray[32][22], dotarray[33][22], dotarray[34][22], dotarray[35][22], dotarray[36][22], dotarray[37][22], dotarray[38][22], dotarray[39][22], dotarray[40][22], dotarray[41][22], dotarray[42][22], dotarray[43][22], dotarray[44][22], dotarray[45][22], dotarray[46][22], dotarray[47][22], dotarray[48][22], dotarray[49][22], dotarray[50][22], dotarray[51][22], dotarray[52][22], dotarray[53][22], dotarray[54][22], dotarray[55][22], dotarray[56][22], dotarray[57][22], dotarray[58][22], dotarray[59][22], dotarray[60][22], dotarray[61][22], dotarray[62][22], dotarray[63][22], dotarray[64][22], dotarray[65][22], dotarray[66][22], dotarray[67][22], dotarray[68][22], dotarray[69][22], dotarray[70][22], dotarray[71][22], dotarray[72][22], dotarray[73][22], dotarray[74][22], dotarray[75][22], dotarray[76][22], dotarray[77][22], dotarray[78][22], dotarray[79][22], dotarray[80][22], dotarray[81][22], dotarray[82][22], dotarray[83][22], dotarray[84][22], dotarray[85][22], dotarray[86][22], dotarray[87][22], dotarray[88][22], dotarray[89][22], dotarray[90][22], dotarray[91][22], dotarray[92][22], dotarray[93][22], dotarray[94][22], dotarray[95][22], dotarray[96][22], dotarray[97][22], dotarray[98][22], dotarray[99][22], dotarray[100][22], dotarray[101][22], dotarray[102][22], dotarray[103][22], dotarray[104][22], dotarray[105][22], dotarray[106][22], dotarray[107][22], dotarray[108][22], dotarray[109][22], dotarray[110][22], dotarray[111][22], dotarray[112][22], dotarray[113][22], dotarray[114][22], dotarray[115][22], dotarray[116][22], dotarray[117][22], dotarray[118][22], dotarray[119][22], dotarray[120][22], dotarray[121][22], dotarray[122][22], dotarray[123][22], dotarray[124][22], dotarray[125][22], dotarray[126][22], dotarray[127][22]};
assign dot_col_23 = {dotarray[0][23], dotarray[1][23], dotarray[2][23], dotarray[3][23], dotarray[4][23], dotarray[5][23], dotarray[6][23], dotarray[7][23], dotarray[8][23], dotarray[9][23], dotarray[10][23], dotarray[11][23], dotarray[12][23], dotarray[13][23], dotarray[14][23], dotarray[15][23], dotarray[16][23], dotarray[17][23], dotarray[18][23], dotarray[19][23], dotarray[20][23], dotarray[21][23], dotarray[22][23], dotarray[23][23], dotarray[24][23], dotarray[25][23], dotarray[26][23], dotarray[27][23], dotarray[28][23], dotarray[29][23], dotarray[30][23], dotarray[31][23], dotarray[32][23], dotarray[33][23], dotarray[34][23], dotarray[35][23], dotarray[36][23], dotarray[37][23], dotarray[38][23], dotarray[39][23], dotarray[40][23], dotarray[41][23], dotarray[42][23], dotarray[43][23], dotarray[44][23], dotarray[45][23], dotarray[46][23], dotarray[47][23], dotarray[48][23], dotarray[49][23], dotarray[50][23], dotarray[51][23], dotarray[52][23], dotarray[53][23], dotarray[54][23], dotarray[55][23], dotarray[56][23], dotarray[57][23], dotarray[58][23], dotarray[59][23], dotarray[60][23], dotarray[61][23], dotarray[62][23], dotarray[63][23], dotarray[64][23], dotarray[65][23], dotarray[66][23], dotarray[67][23], dotarray[68][23], dotarray[69][23], dotarray[70][23], dotarray[71][23], dotarray[72][23], dotarray[73][23], dotarray[74][23], dotarray[75][23], dotarray[76][23], dotarray[77][23], dotarray[78][23], dotarray[79][23], dotarray[80][23], dotarray[81][23], dotarray[82][23], dotarray[83][23], dotarray[84][23], dotarray[85][23], dotarray[86][23], dotarray[87][23], dotarray[88][23], dotarray[89][23], dotarray[90][23], dotarray[91][23], dotarray[92][23], dotarray[93][23], dotarray[94][23], dotarray[95][23], dotarray[96][23], dotarray[97][23], dotarray[98][23], dotarray[99][23], dotarray[100][23], dotarray[101][23], dotarray[102][23], dotarray[103][23], dotarray[104][23], dotarray[105][23], dotarray[106][23], dotarray[107][23], dotarray[108][23], dotarray[109][23], dotarray[110][23], dotarray[111][23], dotarray[112][23], dotarray[113][23], dotarray[114][23], dotarray[115][23], dotarray[116][23], dotarray[117][23], dotarray[118][23], dotarray[119][23], dotarray[120][23], dotarray[121][23], dotarray[122][23], dotarray[123][23], dotarray[124][23], dotarray[125][23], dotarray[126][23], dotarray[127][23]};
assign dot_col_24 = {dotarray[0][24], dotarray[1][24], dotarray[2][24], dotarray[3][24], dotarray[4][24], dotarray[5][24], dotarray[6][24], dotarray[7][24], dotarray[8][24], dotarray[9][24], dotarray[10][24], dotarray[11][24], dotarray[12][24], dotarray[13][24], dotarray[14][24], dotarray[15][24], dotarray[16][24], dotarray[17][24], dotarray[18][24], dotarray[19][24], dotarray[20][24], dotarray[21][24], dotarray[22][24], dotarray[23][24], dotarray[24][24], dotarray[25][24], dotarray[26][24], dotarray[27][24], dotarray[28][24], dotarray[29][24], dotarray[30][24], dotarray[31][24], dotarray[32][24], dotarray[33][24], dotarray[34][24], dotarray[35][24], dotarray[36][24], dotarray[37][24], dotarray[38][24], dotarray[39][24], dotarray[40][24], dotarray[41][24], dotarray[42][24], dotarray[43][24], dotarray[44][24], dotarray[45][24], dotarray[46][24], dotarray[47][24], dotarray[48][24], dotarray[49][24], dotarray[50][24], dotarray[51][24], dotarray[52][24], dotarray[53][24], dotarray[54][24], dotarray[55][24], dotarray[56][24], dotarray[57][24], dotarray[58][24], dotarray[59][24], dotarray[60][24], dotarray[61][24], dotarray[62][24], dotarray[63][24], dotarray[64][24], dotarray[65][24], dotarray[66][24], dotarray[67][24], dotarray[68][24], dotarray[69][24], dotarray[70][24], dotarray[71][24], dotarray[72][24], dotarray[73][24], dotarray[74][24], dotarray[75][24], dotarray[76][24], dotarray[77][24], dotarray[78][24], dotarray[79][24], dotarray[80][24], dotarray[81][24], dotarray[82][24], dotarray[83][24], dotarray[84][24], dotarray[85][24], dotarray[86][24], dotarray[87][24], dotarray[88][24], dotarray[89][24], dotarray[90][24], dotarray[91][24], dotarray[92][24], dotarray[93][24], dotarray[94][24], dotarray[95][24], dotarray[96][24], dotarray[97][24], dotarray[98][24], dotarray[99][24], dotarray[100][24], dotarray[101][24], dotarray[102][24], dotarray[103][24], dotarray[104][24], dotarray[105][24], dotarray[106][24], dotarray[107][24], dotarray[108][24], dotarray[109][24], dotarray[110][24], dotarray[111][24], dotarray[112][24], dotarray[113][24], dotarray[114][24], dotarray[115][24], dotarray[116][24], dotarray[117][24], dotarray[118][24], dotarray[119][24], dotarray[120][24], dotarray[121][24], dotarray[122][24], dotarray[123][24], dotarray[124][24], dotarray[125][24], dotarray[126][24], dotarray[127][24]};
assign dot_col_25 = {dotarray[0][25], dotarray[1][25], dotarray[2][25], dotarray[3][25], dotarray[4][25], dotarray[5][25], dotarray[6][25], dotarray[7][25], dotarray[8][25], dotarray[9][25], dotarray[10][25], dotarray[11][25], dotarray[12][25], dotarray[13][25], dotarray[14][25], dotarray[15][25], dotarray[16][25], dotarray[17][25], dotarray[18][25], dotarray[19][25], dotarray[20][25], dotarray[21][25], dotarray[22][25], dotarray[23][25], dotarray[24][25], dotarray[25][25], dotarray[26][25], dotarray[27][25], dotarray[28][25], dotarray[29][25], dotarray[30][25], dotarray[31][25], dotarray[32][25], dotarray[33][25], dotarray[34][25], dotarray[35][25], dotarray[36][25], dotarray[37][25], dotarray[38][25], dotarray[39][25], dotarray[40][25], dotarray[41][25], dotarray[42][25], dotarray[43][25], dotarray[44][25], dotarray[45][25], dotarray[46][25], dotarray[47][25], dotarray[48][25], dotarray[49][25], dotarray[50][25], dotarray[51][25], dotarray[52][25], dotarray[53][25], dotarray[54][25], dotarray[55][25], dotarray[56][25], dotarray[57][25], dotarray[58][25], dotarray[59][25], dotarray[60][25], dotarray[61][25], dotarray[62][25], dotarray[63][25], dotarray[64][25], dotarray[65][25], dotarray[66][25], dotarray[67][25], dotarray[68][25], dotarray[69][25], dotarray[70][25], dotarray[71][25], dotarray[72][25], dotarray[73][25], dotarray[74][25], dotarray[75][25], dotarray[76][25], dotarray[77][25], dotarray[78][25], dotarray[79][25], dotarray[80][25], dotarray[81][25], dotarray[82][25], dotarray[83][25], dotarray[84][25], dotarray[85][25], dotarray[86][25], dotarray[87][25], dotarray[88][25], dotarray[89][25], dotarray[90][25], dotarray[91][25], dotarray[92][25], dotarray[93][25], dotarray[94][25], dotarray[95][25], dotarray[96][25], dotarray[97][25], dotarray[98][25], dotarray[99][25], dotarray[100][25], dotarray[101][25], dotarray[102][25], dotarray[103][25], dotarray[104][25], dotarray[105][25], dotarray[106][25], dotarray[107][25], dotarray[108][25], dotarray[109][25], dotarray[110][25], dotarray[111][25], dotarray[112][25], dotarray[113][25], dotarray[114][25], dotarray[115][25], dotarray[116][25], dotarray[117][25], dotarray[118][25], dotarray[119][25], dotarray[120][25], dotarray[121][25], dotarray[122][25], dotarray[123][25], dotarray[124][25], dotarray[125][25], dotarray[126][25], dotarray[127][25]};
assign dot_col_26 = {dotarray[0][26], dotarray[1][26], dotarray[2][26], dotarray[3][26], dotarray[4][26], dotarray[5][26], dotarray[6][26], dotarray[7][26], dotarray[8][26], dotarray[9][26], dotarray[10][26], dotarray[11][26], dotarray[12][26], dotarray[13][26], dotarray[14][26], dotarray[15][26], dotarray[16][26], dotarray[17][26], dotarray[18][26], dotarray[19][26], dotarray[20][26], dotarray[21][26], dotarray[22][26], dotarray[23][26], dotarray[24][26], dotarray[25][26], dotarray[26][26], dotarray[27][26], dotarray[28][26], dotarray[29][26], dotarray[30][26], dotarray[31][26], dotarray[32][26], dotarray[33][26], dotarray[34][26], dotarray[35][26], dotarray[36][26], dotarray[37][26], dotarray[38][26], dotarray[39][26], dotarray[40][26], dotarray[41][26], dotarray[42][26], dotarray[43][26], dotarray[44][26], dotarray[45][26], dotarray[46][26], dotarray[47][26], dotarray[48][26], dotarray[49][26], dotarray[50][26], dotarray[51][26], dotarray[52][26], dotarray[53][26], dotarray[54][26], dotarray[55][26], dotarray[56][26], dotarray[57][26], dotarray[58][26], dotarray[59][26], dotarray[60][26], dotarray[61][26], dotarray[62][26], dotarray[63][26], dotarray[64][26], dotarray[65][26], dotarray[66][26], dotarray[67][26], dotarray[68][26], dotarray[69][26], dotarray[70][26], dotarray[71][26], dotarray[72][26], dotarray[73][26], dotarray[74][26], dotarray[75][26], dotarray[76][26], dotarray[77][26], dotarray[78][26], dotarray[79][26], dotarray[80][26], dotarray[81][26], dotarray[82][26], dotarray[83][26], dotarray[84][26], dotarray[85][26], dotarray[86][26], dotarray[87][26], dotarray[88][26], dotarray[89][26], dotarray[90][26], dotarray[91][26], dotarray[92][26], dotarray[93][26], dotarray[94][26], dotarray[95][26], dotarray[96][26], dotarray[97][26], dotarray[98][26], dotarray[99][26], dotarray[100][26], dotarray[101][26], dotarray[102][26], dotarray[103][26], dotarray[104][26], dotarray[105][26], dotarray[106][26], dotarray[107][26], dotarray[108][26], dotarray[109][26], dotarray[110][26], dotarray[111][26], dotarray[112][26], dotarray[113][26], dotarray[114][26], dotarray[115][26], dotarray[116][26], dotarray[117][26], dotarray[118][26], dotarray[119][26], dotarray[120][26], dotarray[121][26], dotarray[122][26], dotarray[123][26], dotarray[124][26], dotarray[125][26], dotarray[126][26], dotarray[127][26]};
assign dot_col_27 = {dotarray[0][27], dotarray[1][27], dotarray[2][27], dotarray[3][27], dotarray[4][27], dotarray[5][27], dotarray[6][27], dotarray[7][27], dotarray[8][27], dotarray[9][27], dotarray[10][27], dotarray[11][27], dotarray[12][27], dotarray[13][27], dotarray[14][27], dotarray[15][27], dotarray[16][27], dotarray[17][27], dotarray[18][27], dotarray[19][27], dotarray[20][27], dotarray[21][27], dotarray[22][27], dotarray[23][27], dotarray[24][27], dotarray[25][27], dotarray[26][27], dotarray[27][27], dotarray[28][27], dotarray[29][27], dotarray[30][27], dotarray[31][27], dotarray[32][27], dotarray[33][27], dotarray[34][27], dotarray[35][27], dotarray[36][27], dotarray[37][27], dotarray[38][27], dotarray[39][27], dotarray[40][27], dotarray[41][27], dotarray[42][27], dotarray[43][27], dotarray[44][27], dotarray[45][27], dotarray[46][27], dotarray[47][27], dotarray[48][27], dotarray[49][27], dotarray[50][27], dotarray[51][27], dotarray[52][27], dotarray[53][27], dotarray[54][27], dotarray[55][27], dotarray[56][27], dotarray[57][27], dotarray[58][27], dotarray[59][27], dotarray[60][27], dotarray[61][27], dotarray[62][27], dotarray[63][27], dotarray[64][27], dotarray[65][27], dotarray[66][27], dotarray[67][27], dotarray[68][27], dotarray[69][27], dotarray[70][27], dotarray[71][27], dotarray[72][27], dotarray[73][27], dotarray[74][27], dotarray[75][27], dotarray[76][27], dotarray[77][27], dotarray[78][27], dotarray[79][27], dotarray[80][27], dotarray[81][27], dotarray[82][27], dotarray[83][27], dotarray[84][27], dotarray[85][27], dotarray[86][27], dotarray[87][27], dotarray[88][27], dotarray[89][27], dotarray[90][27], dotarray[91][27], dotarray[92][27], dotarray[93][27], dotarray[94][27], dotarray[95][27], dotarray[96][27], dotarray[97][27], dotarray[98][27], dotarray[99][27], dotarray[100][27], dotarray[101][27], dotarray[102][27], dotarray[103][27], dotarray[104][27], dotarray[105][27], dotarray[106][27], dotarray[107][27], dotarray[108][27], dotarray[109][27], dotarray[110][27], dotarray[111][27], dotarray[112][27], dotarray[113][27], dotarray[114][27], dotarray[115][27], dotarray[116][27], dotarray[117][27], dotarray[118][27], dotarray[119][27], dotarray[120][27], dotarray[121][27], dotarray[122][27], dotarray[123][27], dotarray[124][27], dotarray[125][27], dotarray[126][27], dotarray[127][27]};
assign dot_col_28 = {dotarray[0][28], dotarray[1][28], dotarray[2][28], dotarray[3][28], dotarray[4][28], dotarray[5][28], dotarray[6][28], dotarray[7][28], dotarray[8][28], dotarray[9][28], dotarray[10][28], dotarray[11][28], dotarray[12][28], dotarray[13][28], dotarray[14][28], dotarray[15][28], dotarray[16][28], dotarray[17][28], dotarray[18][28], dotarray[19][28], dotarray[20][28], dotarray[21][28], dotarray[22][28], dotarray[23][28], dotarray[24][28], dotarray[25][28], dotarray[26][28], dotarray[27][28], dotarray[28][28], dotarray[29][28], dotarray[30][28], dotarray[31][28], dotarray[32][28], dotarray[33][28], dotarray[34][28], dotarray[35][28], dotarray[36][28], dotarray[37][28], dotarray[38][28], dotarray[39][28], dotarray[40][28], dotarray[41][28], dotarray[42][28], dotarray[43][28], dotarray[44][28], dotarray[45][28], dotarray[46][28], dotarray[47][28], dotarray[48][28], dotarray[49][28], dotarray[50][28], dotarray[51][28], dotarray[52][28], dotarray[53][28], dotarray[54][28], dotarray[55][28], dotarray[56][28], dotarray[57][28], dotarray[58][28], dotarray[59][28], dotarray[60][28], dotarray[61][28], dotarray[62][28], dotarray[63][28], dotarray[64][28], dotarray[65][28], dotarray[66][28], dotarray[67][28], dotarray[68][28], dotarray[69][28], dotarray[70][28], dotarray[71][28], dotarray[72][28], dotarray[73][28], dotarray[74][28], dotarray[75][28], dotarray[76][28], dotarray[77][28], dotarray[78][28], dotarray[79][28], dotarray[80][28], dotarray[81][28], dotarray[82][28], dotarray[83][28], dotarray[84][28], dotarray[85][28], dotarray[86][28], dotarray[87][28], dotarray[88][28], dotarray[89][28], dotarray[90][28], dotarray[91][28], dotarray[92][28], dotarray[93][28], dotarray[94][28], dotarray[95][28], dotarray[96][28], dotarray[97][28], dotarray[98][28], dotarray[99][28], dotarray[100][28], dotarray[101][28], dotarray[102][28], dotarray[103][28], dotarray[104][28], dotarray[105][28], dotarray[106][28], dotarray[107][28], dotarray[108][28], dotarray[109][28], dotarray[110][28], dotarray[111][28], dotarray[112][28], dotarray[113][28], dotarray[114][28], dotarray[115][28], dotarray[116][28], dotarray[117][28], dotarray[118][28], dotarray[119][28], dotarray[120][28], dotarray[121][28], dotarray[122][28], dotarray[123][28], dotarray[124][28], dotarray[125][28], dotarray[126][28], dotarray[127][28]};
assign dot_col_29 = {dotarray[0][29], dotarray[1][29], dotarray[2][29], dotarray[3][29], dotarray[4][29], dotarray[5][29], dotarray[6][29], dotarray[7][29], dotarray[8][29], dotarray[9][29], dotarray[10][29], dotarray[11][29], dotarray[12][29], dotarray[13][29], dotarray[14][29], dotarray[15][29], dotarray[16][29], dotarray[17][29], dotarray[18][29], dotarray[19][29], dotarray[20][29], dotarray[21][29], dotarray[22][29], dotarray[23][29], dotarray[24][29], dotarray[25][29], dotarray[26][29], dotarray[27][29], dotarray[28][29], dotarray[29][29], dotarray[30][29], dotarray[31][29], dotarray[32][29], dotarray[33][29], dotarray[34][29], dotarray[35][29], dotarray[36][29], dotarray[37][29], dotarray[38][29], dotarray[39][29], dotarray[40][29], dotarray[41][29], dotarray[42][29], dotarray[43][29], dotarray[44][29], dotarray[45][29], dotarray[46][29], dotarray[47][29], dotarray[48][29], dotarray[49][29], dotarray[50][29], dotarray[51][29], dotarray[52][29], dotarray[53][29], dotarray[54][29], dotarray[55][29], dotarray[56][29], dotarray[57][29], dotarray[58][29], dotarray[59][29], dotarray[60][29], dotarray[61][29], dotarray[62][29], dotarray[63][29], dotarray[64][29], dotarray[65][29], dotarray[66][29], dotarray[67][29], dotarray[68][29], dotarray[69][29], dotarray[70][29], dotarray[71][29], dotarray[72][29], dotarray[73][29], dotarray[74][29], dotarray[75][29], dotarray[76][29], dotarray[77][29], dotarray[78][29], dotarray[79][29], dotarray[80][29], dotarray[81][29], dotarray[82][29], dotarray[83][29], dotarray[84][29], dotarray[85][29], dotarray[86][29], dotarray[87][29], dotarray[88][29], dotarray[89][29], dotarray[90][29], dotarray[91][29], dotarray[92][29], dotarray[93][29], dotarray[94][29], dotarray[95][29], dotarray[96][29], dotarray[97][29], dotarray[98][29], dotarray[99][29], dotarray[100][29], dotarray[101][29], dotarray[102][29], dotarray[103][29], dotarray[104][29], dotarray[105][29], dotarray[106][29], dotarray[107][29], dotarray[108][29], dotarray[109][29], dotarray[110][29], dotarray[111][29], dotarray[112][29], dotarray[113][29], dotarray[114][29], dotarray[115][29], dotarray[116][29], dotarray[117][29], dotarray[118][29], dotarray[119][29], dotarray[120][29], dotarray[121][29], dotarray[122][29], dotarray[123][29], dotarray[124][29], dotarray[125][29], dotarray[126][29], dotarray[127][29]};
assign dot_col_30 = {dotarray[0][30], dotarray[1][30], dotarray[2][30], dotarray[3][30], dotarray[4][30], dotarray[5][30], dotarray[6][30], dotarray[7][30], dotarray[8][30], dotarray[9][30], dotarray[10][30], dotarray[11][30], dotarray[12][30], dotarray[13][30], dotarray[14][30], dotarray[15][30], dotarray[16][30], dotarray[17][30], dotarray[18][30], dotarray[19][30], dotarray[20][30], dotarray[21][30], dotarray[22][30], dotarray[23][30], dotarray[24][30], dotarray[25][30], dotarray[26][30], dotarray[27][30], dotarray[28][30], dotarray[29][30], dotarray[30][30], dotarray[31][30], dotarray[32][30], dotarray[33][30], dotarray[34][30], dotarray[35][30], dotarray[36][30], dotarray[37][30], dotarray[38][30], dotarray[39][30], dotarray[40][30], dotarray[41][30], dotarray[42][30], dotarray[43][30], dotarray[44][30], dotarray[45][30], dotarray[46][30], dotarray[47][30], dotarray[48][30], dotarray[49][30], dotarray[50][30], dotarray[51][30], dotarray[52][30], dotarray[53][30], dotarray[54][30], dotarray[55][30], dotarray[56][30], dotarray[57][30], dotarray[58][30], dotarray[59][30], dotarray[60][30], dotarray[61][30], dotarray[62][30], dotarray[63][30], dotarray[64][30], dotarray[65][30], dotarray[66][30], dotarray[67][30], dotarray[68][30], dotarray[69][30], dotarray[70][30], dotarray[71][30], dotarray[72][30], dotarray[73][30], dotarray[74][30], dotarray[75][30], dotarray[76][30], dotarray[77][30], dotarray[78][30], dotarray[79][30], dotarray[80][30], dotarray[81][30], dotarray[82][30], dotarray[83][30], dotarray[84][30], dotarray[85][30], dotarray[86][30], dotarray[87][30], dotarray[88][30], dotarray[89][30], dotarray[90][30], dotarray[91][30], dotarray[92][30], dotarray[93][30], dotarray[94][30], dotarray[95][30], dotarray[96][30], dotarray[97][30], dotarray[98][30], dotarray[99][30], dotarray[100][30], dotarray[101][30], dotarray[102][30], dotarray[103][30], dotarray[104][30], dotarray[105][30], dotarray[106][30], dotarray[107][30], dotarray[108][30], dotarray[109][30], dotarray[110][30], dotarray[111][30], dotarray[112][30], dotarray[113][30], dotarray[114][30], dotarray[115][30], dotarray[116][30], dotarray[117][30], dotarray[118][30], dotarray[119][30], dotarray[120][30], dotarray[121][30], dotarray[122][30], dotarray[123][30], dotarray[124][30], dotarray[125][30], dotarray[126][30], dotarray[127][30]};
assign dot_col_31 = {dotarray[0][31], dotarray[1][31], dotarray[2][31], dotarray[3][31], dotarray[4][31], dotarray[5][31], dotarray[6][31], dotarray[7][31], dotarray[8][31], dotarray[9][31], dotarray[10][31], dotarray[11][31], dotarray[12][31], dotarray[13][31], dotarray[14][31], dotarray[15][31], dotarray[16][31], dotarray[17][31], dotarray[18][31], dotarray[19][31], dotarray[20][31], dotarray[21][31], dotarray[22][31], dotarray[23][31], dotarray[24][31], dotarray[25][31], dotarray[26][31], dotarray[27][31], dotarray[28][31], dotarray[29][31], dotarray[30][31], dotarray[31][31], dotarray[32][31], dotarray[33][31], dotarray[34][31], dotarray[35][31], dotarray[36][31], dotarray[37][31], dotarray[38][31], dotarray[39][31], dotarray[40][31], dotarray[41][31], dotarray[42][31], dotarray[43][31], dotarray[44][31], dotarray[45][31], dotarray[46][31], dotarray[47][31], dotarray[48][31], dotarray[49][31], dotarray[50][31], dotarray[51][31], dotarray[52][31], dotarray[53][31], dotarray[54][31], dotarray[55][31], dotarray[56][31], dotarray[57][31], dotarray[58][31], dotarray[59][31], dotarray[60][31], dotarray[61][31], dotarray[62][31], dotarray[63][31], dotarray[64][31], dotarray[65][31], dotarray[66][31], dotarray[67][31], dotarray[68][31], dotarray[69][31], dotarray[70][31], dotarray[71][31], dotarray[72][31], dotarray[73][31], dotarray[74][31], dotarray[75][31], dotarray[76][31], dotarray[77][31], dotarray[78][31], dotarray[79][31], dotarray[80][31], dotarray[81][31], dotarray[82][31], dotarray[83][31], dotarray[84][31], dotarray[85][31], dotarray[86][31], dotarray[87][31], dotarray[88][31], dotarray[89][31], dotarray[90][31], dotarray[91][31], dotarray[92][31], dotarray[93][31], dotarray[94][31], dotarray[95][31], dotarray[96][31], dotarray[97][31], dotarray[98][31], dotarray[99][31], dotarray[100][31], dotarray[101][31], dotarray[102][31], dotarray[103][31], dotarray[104][31], dotarray[105][31], dotarray[106][31], dotarray[107][31], dotarray[108][31], dotarray[109][31], dotarray[110][31], dotarray[111][31], dotarray[112][31], dotarray[113][31], dotarray[114][31], dotarray[115][31], dotarray[116][31], dotarray[117][31], dotarray[118][31], dotarray[119][31], dotarray[120][31], dotarray[121][31], dotarray[122][31], dotarray[123][31], dotarray[124][31], dotarray[125][31], dotarray[126][31], dotarray[127][31]};
assign dot_col_32 = {dotarray[0][32], dotarray[1][32], dotarray[2][32], dotarray[3][32], dotarray[4][32], dotarray[5][32], dotarray[6][32], dotarray[7][32], dotarray[8][32], dotarray[9][32], dotarray[10][32], dotarray[11][32], dotarray[12][32], dotarray[13][32], dotarray[14][32], dotarray[15][32], dotarray[16][32], dotarray[17][32], dotarray[18][32], dotarray[19][32], dotarray[20][32], dotarray[21][32], dotarray[22][32], dotarray[23][32], dotarray[24][32], dotarray[25][32], dotarray[26][32], dotarray[27][32], dotarray[28][32], dotarray[29][32], dotarray[30][32], dotarray[31][32], dotarray[32][32], dotarray[33][32], dotarray[34][32], dotarray[35][32], dotarray[36][32], dotarray[37][32], dotarray[38][32], dotarray[39][32], dotarray[40][32], dotarray[41][32], dotarray[42][32], dotarray[43][32], dotarray[44][32], dotarray[45][32], dotarray[46][32], dotarray[47][32], dotarray[48][32], dotarray[49][32], dotarray[50][32], dotarray[51][32], dotarray[52][32], dotarray[53][32], dotarray[54][32], dotarray[55][32], dotarray[56][32], dotarray[57][32], dotarray[58][32], dotarray[59][32], dotarray[60][32], dotarray[61][32], dotarray[62][32], dotarray[63][32], dotarray[64][32], dotarray[65][32], dotarray[66][32], dotarray[67][32], dotarray[68][32], dotarray[69][32], dotarray[70][32], dotarray[71][32], dotarray[72][32], dotarray[73][32], dotarray[74][32], dotarray[75][32], dotarray[76][32], dotarray[77][32], dotarray[78][32], dotarray[79][32], dotarray[80][32], dotarray[81][32], dotarray[82][32], dotarray[83][32], dotarray[84][32], dotarray[85][32], dotarray[86][32], dotarray[87][32], dotarray[88][32], dotarray[89][32], dotarray[90][32], dotarray[91][32], dotarray[92][32], dotarray[93][32], dotarray[94][32], dotarray[95][32], dotarray[96][32], dotarray[97][32], dotarray[98][32], dotarray[99][32], dotarray[100][32], dotarray[101][32], dotarray[102][32], dotarray[103][32], dotarray[104][32], dotarray[105][32], dotarray[106][32], dotarray[107][32], dotarray[108][32], dotarray[109][32], dotarray[110][32], dotarray[111][32], dotarray[112][32], dotarray[113][32], dotarray[114][32], dotarray[115][32], dotarray[116][32], dotarray[117][32], dotarray[118][32], dotarray[119][32], dotarray[120][32], dotarray[121][32], dotarray[122][32], dotarray[123][32], dotarray[124][32], dotarray[125][32], dotarray[126][32], dotarray[127][32]};
assign dot_col_33 = {dotarray[0][33], dotarray[1][33], dotarray[2][33], dotarray[3][33], dotarray[4][33], dotarray[5][33], dotarray[6][33], dotarray[7][33], dotarray[8][33], dotarray[9][33], dotarray[10][33], dotarray[11][33], dotarray[12][33], dotarray[13][33], dotarray[14][33], dotarray[15][33], dotarray[16][33], dotarray[17][33], dotarray[18][33], dotarray[19][33], dotarray[20][33], dotarray[21][33], dotarray[22][33], dotarray[23][33], dotarray[24][33], dotarray[25][33], dotarray[26][33], dotarray[27][33], dotarray[28][33], dotarray[29][33], dotarray[30][33], dotarray[31][33], dotarray[32][33], dotarray[33][33], dotarray[34][33], dotarray[35][33], dotarray[36][33], dotarray[37][33], dotarray[38][33], dotarray[39][33], dotarray[40][33], dotarray[41][33], dotarray[42][33], dotarray[43][33], dotarray[44][33], dotarray[45][33], dotarray[46][33], dotarray[47][33], dotarray[48][33], dotarray[49][33], dotarray[50][33], dotarray[51][33], dotarray[52][33], dotarray[53][33], dotarray[54][33], dotarray[55][33], dotarray[56][33], dotarray[57][33], dotarray[58][33], dotarray[59][33], dotarray[60][33], dotarray[61][33], dotarray[62][33], dotarray[63][33], dotarray[64][33], dotarray[65][33], dotarray[66][33], dotarray[67][33], dotarray[68][33], dotarray[69][33], dotarray[70][33], dotarray[71][33], dotarray[72][33], dotarray[73][33], dotarray[74][33], dotarray[75][33], dotarray[76][33], dotarray[77][33], dotarray[78][33], dotarray[79][33], dotarray[80][33], dotarray[81][33], dotarray[82][33], dotarray[83][33], dotarray[84][33], dotarray[85][33], dotarray[86][33], dotarray[87][33], dotarray[88][33], dotarray[89][33], dotarray[90][33], dotarray[91][33], dotarray[92][33], dotarray[93][33], dotarray[94][33], dotarray[95][33], dotarray[96][33], dotarray[97][33], dotarray[98][33], dotarray[99][33], dotarray[100][33], dotarray[101][33], dotarray[102][33], dotarray[103][33], dotarray[104][33], dotarray[105][33], dotarray[106][33], dotarray[107][33], dotarray[108][33], dotarray[109][33], dotarray[110][33], dotarray[111][33], dotarray[112][33], dotarray[113][33], dotarray[114][33], dotarray[115][33], dotarray[116][33], dotarray[117][33], dotarray[118][33], dotarray[119][33], dotarray[120][33], dotarray[121][33], dotarray[122][33], dotarray[123][33], dotarray[124][33], dotarray[125][33], dotarray[126][33], dotarray[127][33]};
assign dot_col_34 = {dotarray[0][34], dotarray[1][34], dotarray[2][34], dotarray[3][34], dotarray[4][34], dotarray[5][34], dotarray[6][34], dotarray[7][34], dotarray[8][34], dotarray[9][34], dotarray[10][34], dotarray[11][34], dotarray[12][34], dotarray[13][34], dotarray[14][34], dotarray[15][34], dotarray[16][34], dotarray[17][34], dotarray[18][34], dotarray[19][34], dotarray[20][34], dotarray[21][34], dotarray[22][34], dotarray[23][34], dotarray[24][34], dotarray[25][34], dotarray[26][34], dotarray[27][34], dotarray[28][34], dotarray[29][34], dotarray[30][34], dotarray[31][34], dotarray[32][34], dotarray[33][34], dotarray[34][34], dotarray[35][34], dotarray[36][34], dotarray[37][34], dotarray[38][34], dotarray[39][34], dotarray[40][34], dotarray[41][34], dotarray[42][34], dotarray[43][34], dotarray[44][34], dotarray[45][34], dotarray[46][34], dotarray[47][34], dotarray[48][34], dotarray[49][34], dotarray[50][34], dotarray[51][34], dotarray[52][34], dotarray[53][34], dotarray[54][34], dotarray[55][34], dotarray[56][34], dotarray[57][34], dotarray[58][34], dotarray[59][34], dotarray[60][34], dotarray[61][34], dotarray[62][34], dotarray[63][34], dotarray[64][34], dotarray[65][34], dotarray[66][34], dotarray[67][34], dotarray[68][34], dotarray[69][34], dotarray[70][34], dotarray[71][34], dotarray[72][34], dotarray[73][34], dotarray[74][34], dotarray[75][34], dotarray[76][34], dotarray[77][34], dotarray[78][34], dotarray[79][34], dotarray[80][34], dotarray[81][34], dotarray[82][34], dotarray[83][34], dotarray[84][34], dotarray[85][34], dotarray[86][34], dotarray[87][34], dotarray[88][34], dotarray[89][34], dotarray[90][34], dotarray[91][34], dotarray[92][34], dotarray[93][34], dotarray[94][34], dotarray[95][34], dotarray[96][34], dotarray[97][34], dotarray[98][34], dotarray[99][34], dotarray[100][34], dotarray[101][34], dotarray[102][34], dotarray[103][34], dotarray[104][34], dotarray[105][34], dotarray[106][34], dotarray[107][34], dotarray[108][34], dotarray[109][34], dotarray[110][34], dotarray[111][34], dotarray[112][34], dotarray[113][34], dotarray[114][34], dotarray[115][34], dotarray[116][34], dotarray[117][34], dotarray[118][34], dotarray[119][34], dotarray[120][34], dotarray[121][34], dotarray[122][34], dotarray[123][34], dotarray[124][34], dotarray[125][34], dotarray[126][34], dotarray[127][34]};
assign dot_col_35 = {dotarray[0][35], dotarray[1][35], dotarray[2][35], dotarray[3][35], dotarray[4][35], dotarray[5][35], dotarray[6][35], dotarray[7][35], dotarray[8][35], dotarray[9][35], dotarray[10][35], dotarray[11][35], dotarray[12][35], dotarray[13][35], dotarray[14][35], dotarray[15][35], dotarray[16][35], dotarray[17][35], dotarray[18][35], dotarray[19][35], dotarray[20][35], dotarray[21][35], dotarray[22][35], dotarray[23][35], dotarray[24][35], dotarray[25][35], dotarray[26][35], dotarray[27][35], dotarray[28][35], dotarray[29][35], dotarray[30][35], dotarray[31][35], dotarray[32][35], dotarray[33][35], dotarray[34][35], dotarray[35][35], dotarray[36][35], dotarray[37][35], dotarray[38][35], dotarray[39][35], dotarray[40][35], dotarray[41][35], dotarray[42][35], dotarray[43][35], dotarray[44][35], dotarray[45][35], dotarray[46][35], dotarray[47][35], dotarray[48][35], dotarray[49][35], dotarray[50][35], dotarray[51][35], dotarray[52][35], dotarray[53][35], dotarray[54][35], dotarray[55][35], dotarray[56][35], dotarray[57][35], dotarray[58][35], dotarray[59][35], dotarray[60][35], dotarray[61][35], dotarray[62][35], dotarray[63][35], dotarray[64][35], dotarray[65][35], dotarray[66][35], dotarray[67][35], dotarray[68][35], dotarray[69][35], dotarray[70][35], dotarray[71][35], dotarray[72][35], dotarray[73][35], dotarray[74][35], dotarray[75][35], dotarray[76][35], dotarray[77][35], dotarray[78][35], dotarray[79][35], dotarray[80][35], dotarray[81][35], dotarray[82][35], dotarray[83][35], dotarray[84][35], dotarray[85][35], dotarray[86][35], dotarray[87][35], dotarray[88][35], dotarray[89][35], dotarray[90][35], dotarray[91][35], dotarray[92][35], dotarray[93][35], dotarray[94][35], dotarray[95][35], dotarray[96][35], dotarray[97][35], dotarray[98][35], dotarray[99][35], dotarray[100][35], dotarray[101][35], dotarray[102][35], dotarray[103][35], dotarray[104][35], dotarray[105][35], dotarray[106][35], dotarray[107][35], dotarray[108][35], dotarray[109][35], dotarray[110][35], dotarray[111][35], dotarray[112][35], dotarray[113][35], dotarray[114][35], dotarray[115][35], dotarray[116][35], dotarray[117][35], dotarray[118][35], dotarray[119][35], dotarray[120][35], dotarray[121][35], dotarray[122][35], dotarray[123][35], dotarray[124][35], dotarray[125][35], dotarray[126][35], dotarray[127][35]};
assign dot_col_36 = {dotarray[0][36], dotarray[1][36], dotarray[2][36], dotarray[3][36], dotarray[4][36], dotarray[5][36], dotarray[6][36], dotarray[7][36], dotarray[8][36], dotarray[9][36], dotarray[10][36], dotarray[11][36], dotarray[12][36], dotarray[13][36], dotarray[14][36], dotarray[15][36], dotarray[16][36], dotarray[17][36], dotarray[18][36], dotarray[19][36], dotarray[20][36], dotarray[21][36], dotarray[22][36], dotarray[23][36], dotarray[24][36], dotarray[25][36], dotarray[26][36], dotarray[27][36], dotarray[28][36], dotarray[29][36], dotarray[30][36], dotarray[31][36], dotarray[32][36], dotarray[33][36], dotarray[34][36], dotarray[35][36], dotarray[36][36], dotarray[37][36], dotarray[38][36], dotarray[39][36], dotarray[40][36], dotarray[41][36], dotarray[42][36], dotarray[43][36], dotarray[44][36], dotarray[45][36], dotarray[46][36], dotarray[47][36], dotarray[48][36], dotarray[49][36], dotarray[50][36], dotarray[51][36], dotarray[52][36], dotarray[53][36], dotarray[54][36], dotarray[55][36], dotarray[56][36], dotarray[57][36], dotarray[58][36], dotarray[59][36], dotarray[60][36], dotarray[61][36], dotarray[62][36], dotarray[63][36], dotarray[64][36], dotarray[65][36], dotarray[66][36], dotarray[67][36], dotarray[68][36], dotarray[69][36], dotarray[70][36], dotarray[71][36], dotarray[72][36], dotarray[73][36], dotarray[74][36], dotarray[75][36], dotarray[76][36], dotarray[77][36], dotarray[78][36], dotarray[79][36], dotarray[80][36], dotarray[81][36], dotarray[82][36], dotarray[83][36], dotarray[84][36], dotarray[85][36], dotarray[86][36], dotarray[87][36], dotarray[88][36], dotarray[89][36], dotarray[90][36], dotarray[91][36], dotarray[92][36], dotarray[93][36], dotarray[94][36], dotarray[95][36], dotarray[96][36], dotarray[97][36], dotarray[98][36], dotarray[99][36], dotarray[100][36], dotarray[101][36], dotarray[102][36], dotarray[103][36], dotarray[104][36], dotarray[105][36], dotarray[106][36], dotarray[107][36], dotarray[108][36], dotarray[109][36], dotarray[110][36], dotarray[111][36], dotarray[112][36], dotarray[113][36], dotarray[114][36], dotarray[115][36], dotarray[116][36], dotarray[117][36], dotarray[118][36], dotarray[119][36], dotarray[120][36], dotarray[121][36], dotarray[122][36], dotarray[123][36], dotarray[124][36], dotarray[125][36], dotarray[126][36], dotarray[127][36]};
assign dot_col_37 = {dotarray[0][37], dotarray[1][37], dotarray[2][37], dotarray[3][37], dotarray[4][37], dotarray[5][37], dotarray[6][37], dotarray[7][37], dotarray[8][37], dotarray[9][37], dotarray[10][37], dotarray[11][37], dotarray[12][37], dotarray[13][37], dotarray[14][37], dotarray[15][37], dotarray[16][37], dotarray[17][37], dotarray[18][37], dotarray[19][37], dotarray[20][37], dotarray[21][37], dotarray[22][37], dotarray[23][37], dotarray[24][37], dotarray[25][37], dotarray[26][37], dotarray[27][37], dotarray[28][37], dotarray[29][37], dotarray[30][37], dotarray[31][37], dotarray[32][37], dotarray[33][37], dotarray[34][37], dotarray[35][37], dotarray[36][37], dotarray[37][37], dotarray[38][37], dotarray[39][37], dotarray[40][37], dotarray[41][37], dotarray[42][37], dotarray[43][37], dotarray[44][37], dotarray[45][37], dotarray[46][37], dotarray[47][37], dotarray[48][37], dotarray[49][37], dotarray[50][37], dotarray[51][37], dotarray[52][37], dotarray[53][37], dotarray[54][37], dotarray[55][37], dotarray[56][37], dotarray[57][37], dotarray[58][37], dotarray[59][37], dotarray[60][37], dotarray[61][37], dotarray[62][37], dotarray[63][37], dotarray[64][37], dotarray[65][37], dotarray[66][37], dotarray[67][37], dotarray[68][37], dotarray[69][37], dotarray[70][37], dotarray[71][37], dotarray[72][37], dotarray[73][37], dotarray[74][37], dotarray[75][37], dotarray[76][37], dotarray[77][37], dotarray[78][37], dotarray[79][37], dotarray[80][37], dotarray[81][37], dotarray[82][37], dotarray[83][37], dotarray[84][37], dotarray[85][37], dotarray[86][37], dotarray[87][37], dotarray[88][37], dotarray[89][37], dotarray[90][37], dotarray[91][37], dotarray[92][37], dotarray[93][37], dotarray[94][37], dotarray[95][37], dotarray[96][37], dotarray[97][37], dotarray[98][37], dotarray[99][37], dotarray[100][37], dotarray[101][37], dotarray[102][37], dotarray[103][37], dotarray[104][37], dotarray[105][37], dotarray[106][37], dotarray[107][37], dotarray[108][37], dotarray[109][37], dotarray[110][37], dotarray[111][37], dotarray[112][37], dotarray[113][37], dotarray[114][37], dotarray[115][37], dotarray[116][37], dotarray[117][37], dotarray[118][37], dotarray[119][37], dotarray[120][37], dotarray[121][37], dotarray[122][37], dotarray[123][37], dotarray[124][37], dotarray[125][37], dotarray[126][37], dotarray[127][37]};
assign dot_col_38 = {dotarray[0][38], dotarray[1][38], dotarray[2][38], dotarray[3][38], dotarray[4][38], dotarray[5][38], dotarray[6][38], dotarray[7][38], dotarray[8][38], dotarray[9][38], dotarray[10][38], dotarray[11][38], dotarray[12][38], dotarray[13][38], dotarray[14][38], dotarray[15][38], dotarray[16][38], dotarray[17][38], dotarray[18][38], dotarray[19][38], dotarray[20][38], dotarray[21][38], dotarray[22][38], dotarray[23][38], dotarray[24][38], dotarray[25][38], dotarray[26][38], dotarray[27][38], dotarray[28][38], dotarray[29][38], dotarray[30][38], dotarray[31][38], dotarray[32][38], dotarray[33][38], dotarray[34][38], dotarray[35][38], dotarray[36][38], dotarray[37][38], dotarray[38][38], dotarray[39][38], dotarray[40][38], dotarray[41][38], dotarray[42][38], dotarray[43][38], dotarray[44][38], dotarray[45][38], dotarray[46][38], dotarray[47][38], dotarray[48][38], dotarray[49][38], dotarray[50][38], dotarray[51][38], dotarray[52][38], dotarray[53][38], dotarray[54][38], dotarray[55][38], dotarray[56][38], dotarray[57][38], dotarray[58][38], dotarray[59][38], dotarray[60][38], dotarray[61][38], dotarray[62][38], dotarray[63][38], dotarray[64][38], dotarray[65][38], dotarray[66][38], dotarray[67][38], dotarray[68][38], dotarray[69][38], dotarray[70][38], dotarray[71][38], dotarray[72][38], dotarray[73][38], dotarray[74][38], dotarray[75][38], dotarray[76][38], dotarray[77][38], dotarray[78][38], dotarray[79][38], dotarray[80][38], dotarray[81][38], dotarray[82][38], dotarray[83][38], dotarray[84][38], dotarray[85][38], dotarray[86][38], dotarray[87][38], dotarray[88][38], dotarray[89][38], dotarray[90][38], dotarray[91][38], dotarray[92][38], dotarray[93][38], dotarray[94][38], dotarray[95][38], dotarray[96][38], dotarray[97][38], dotarray[98][38], dotarray[99][38], dotarray[100][38], dotarray[101][38], dotarray[102][38], dotarray[103][38], dotarray[104][38], dotarray[105][38], dotarray[106][38], dotarray[107][38], dotarray[108][38], dotarray[109][38], dotarray[110][38], dotarray[111][38], dotarray[112][38], dotarray[113][38], dotarray[114][38], dotarray[115][38], dotarray[116][38], dotarray[117][38], dotarray[118][38], dotarray[119][38], dotarray[120][38], dotarray[121][38], dotarray[122][38], dotarray[123][38], dotarray[124][38], dotarray[125][38], dotarray[126][38], dotarray[127][38]};
assign dot_col_39 = {dotarray[0][39], dotarray[1][39], dotarray[2][39], dotarray[3][39], dotarray[4][39], dotarray[5][39], dotarray[6][39], dotarray[7][39], dotarray[8][39], dotarray[9][39], dotarray[10][39], dotarray[11][39], dotarray[12][39], dotarray[13][39], dotarray[14][39], dotarray[15][39], dotarray[16][39], dotarray[17][39], dotarray[18][39], dotarray[19][39], dotarray[20][39], dotarray[21][39], dotarray[22][39], dotarray[23][39], dotarray[24][39], dotarray[25][39], dotarray[26][39], dotarray[27][39], dotarray[28][39], dotarray[29][39], dotarray[30][39], dotarray[31][39], dotarray[32][39], dotarray[33][39], dotarray[34][39], dotarray[35][39], dotarray[36][39], dotarray[37][39], dotarray[38][39], dotarray[39][39], dotarray[40][39], dotarray[41][39], dotarray[42][39], dotarray[43][39], dotarray[44][39], dotarray[45][39], dotarray[46][39], dotarray[47][39], dotarray[48][39], dotarray[49][39], dotarray[50][39], dotarray[51][39], dotarray[52][39], dotarray[53][39], dotarray[54][39], dotarray[55][39], dotarray[56][39], dotarray[57][39], dotarray[58][39], dotarray[59][39], dotarray[60][39], dotarray[61][39], dotarray[62][39], dotarray[63][39], dotarray[64][39], dotarray[65][39], dotarray[66][39], dotarray[67][39], dotarray[68][39], dotarray[69][39], dotarray[70][39], dotarray[71][39], dotarray[72][39], dotarray[73][39], dotarray[74][39], dotarray[75][39], dotarray[76][39], dotarray[77][39], dotarray[78][39], dotarray[79][39], dotarray[80][39], dotarray[81][39], dotarray[82][39], dotarray[83][39], dotarray[84][39], dotarray[85][39], dotarray[86][39], dotarray[87][39], dotarray[88][39], dotarray[89][39], dotarray[90][39], dotarray[91][39], dotarray[92][39], dotarray[93][39], dotarray[94][39], dotarray[95][39], dotarray[96][39], dotarray[97][39], dotarray[98][39], dotarray[99][39], dotarray[100][39], dotarray[101][39], dotarray[102][39], dotarray[103][39], dotarray[104][39], dotarray[105][39], dotarray[106][39], dotarray[107][39], dotarray[108][39], dotarray[109][39], dotarray[110][39], dotarray[111][39], dotarray[112][39], dotarray[113][39], dotarray[114][39], dotarray[115][39], dotarray[116][39], dotarray[117][39], dotarray[118][39], dotarray[119][39], dotarray[120][39], dotarray[121][39], dotarray[122][39], dotarray[123][39], dotarray[124][39], dotarray[125][39], dotarray[126][39], dotarray[127][39]};
assign dot_col_40 = {dotarray[0][40], dotarray[1][40], dotarray[2][40], dotarray[3][40], dotarray[4][40], dotarray[5][40], dotarray[6][40], dotarray[7][40], dotarray[8][40], dotarray[9][40], dotarray[10][40], dotarray[11][40], dotarray[12][40], dotarray[13][40], dotarray[14][40], dotarray[15][40], dotarray[16][40], dotarray[17][40], dotarray[18][40], dotarray[19][40], dotarray[20][40], dotarray[21][40], dotarray[22][40], dotarray[23][40], dotarray[24][40], dotarray[25][40], dotarray[26][40], dotarray[27][40], dotarray[28][40], dotarray[29][40], dotarray[30][40], dotarray[31][40], dotarray[32][40], dotarray[33][40], dotarray[34][40], dotarray[35][40], dotarray[36][40], dotarray[37][40], dotarray[38][40], dotarray[39][40], dotarray[40][40], dotarray[41][40], dotarray[42][40], dotarray[43][40], dotarray[44][40], dotarray[45][40], dotarray[46][40], dotarray[47][40], dotarray[48][40], dotarray[49][40], dotarray[50][40], dotarray[51][40], dotarray[52][40], dotarray[53][40], dotarray[54][40], dotarray[55][40], dotarray[56][40], dotarray[57][40], dotarray[58][40], dotarray[59][40], dotarray[60][40], dotarray[61][40], dotarray[62][40], dotarray[63][40], dotarray[64][40], dotarray[65][40], dotarray[66][40], dotarray[67][40], dotarray[68][40], dotarray[69][40], dotarray[70][40], dotarray[71][40], dotarray[72][40], dotarray[73][40], dotarray[74][40], dotarray[75][40], dotarray[76][40], dotarray[77][40], dotarray[78][40], dotarray[79][40], dotarray[80][40], dotarray[81][40], dotarray[82][40], dotarray[83][40], dotarray[84][40], dotarray[85][40], dotarray[86][40], dotarray[87][40], dotarray[88][40], dotarray[89][40], dotarray[90][40], dotarray[91][40], dotarray[92][40], dotarray[93][40], dotarray[94][40], dotarray[95][40], dotarray[96][40], dotarray[97][40], dotarray[98][40], dotarray[99][40], dotarray[100][40], dotarray[101][40], dotarray[102][40], dotarray[103][40], dotarray[104][40], dotarray[105][40], dotarray[106][40], dotarray[107][40], dotarray[108][40], dotarray[109][40], dotarray[110][40], dotarray[111][40], dotarray[112][40], dotarray[113][40], dotarray[114][40], dotarray[115][40], dotarray[116][40], dotarray[117][40], dotarray[118][40], dotarray[119][40], dotarray[120][40], dotarray[121][40], dotarray[122][40], dotarray[123][40], dotarray[124][40], dotarray[125][40], dotarray[126][40], dotarray[127][40]};
assign dot_col_41 = {dotarray[0][41], dotarray[1][41], dotarray[2][41], dotarray[3][41], dotarray[4][41], dotarray[5][41], dotarray[6][41], dotarray[7][41], dotarray[8][41], dotarray[9][41], dotarray[10][41], dotarray[11][41], dotarray[12][41], dotarray[13][41], dotarray[14][41], dotarray[15][41], dotarray[16][41], dotarray[17][41], dotarray[18][41], dotarray[19][41], dotarray[20][41], dotarray[21][41], dotarray[22][41], dotarray[23][41], dotarray[24][41], dotarray[25][41], dotarray[26][41], dotarray[27][41], dotarray[28][41], dotarray[29][41], dotarray[30][41], dotarray[31][41], dotarray[32][41], dotarray[33][41], dotarray[34][41], dotarray[35][41], dotarray[36][41], dotarray[37][41], dotarray[38][41], dotarray[39][41], dotarray[40][41], dotarray[41][41], dotarray[42][41], dotarray[43][41], dotarray[44][41], dotarray[45][41], dotarray[46][41], dotarray[47][41], dotarray[48][41], dotarray[49][41], dotarray[50][41], dotarray[51][41], dotarray[52][41], dotarray[53][41], dotarray[54][41], dotarray[55][41], dotarray[56][41], dotarray[57][41], dotarray[58][41], dotarray[59][41], dotarray[60][41], dotarray[61][41], dotarray[62][41], dotarray[63][41], dotarray[64][41], dotarray[65][41], dotarray[66][41], dotarray[67][41], dotarray[68][41], dotarray[69][41], dotarray[70][41], dotarray[71][41], dotarray[72][41], dotarray[73][41], dotarray[74][41], dotarray[75][41], dotarray[76][41], dotarray[77][41], dotarray[78][41], dotarray[79][41], dotarray[80][41], dotarray[81][41], dotarray[82][41], dotarray[83][41], dotarray[84][41], dotarray[85][41], dotarray[86][41], dotarray[87][41], dotarray[88][41], dotarray[89][41], dotarray[90][41], dotarray[91][41], dotarray[92][41], dotarray[93][41], dotarray[94][41], dotarray[95][41], dotarray[96][41], dotarray[97][41], dotarray[98][41], dotarray[99][41], dotarray[100][41], dotarray[101][41], dotarray[102][41], dotarray[103][41], dotarray[104][41], dotarray[105][41], dotarray[106][41], dotarray[107][41], dotarray[108][41], dotarray[109][41], dotarray[110][41], dotarray[111][41], dotarray[112][41], dotarray[113][41], dotarray[114][41], dotarray[115][41], dotarray[116][41], dotarray[117][41], dotarray[118][41], dotarray[119][41], dotarray[120][41], dotarray[121][41], dotarray[122][41], dotarray[123][41], dotarray[124][41], dotarray[125][41], dotarray[126][41], dotarray[127][41]};
assign dot_col_42 = {dotarray[0][42], dotarray[1][42], dotarray[2][42], dotarray[3][42], dotarray[4][42], dotarray[5][42], dotarray[6][42], dotarray[7][42], dotarray[8][42], dotarray[9][42], dotarray[10][42], dotarray[11][42], dotarray[12][42], dotarray[13][42], dotarray[14][42], dotarray[15][42], dotarray[16][42], dotarray[17][42], dotarray[18][42], dotarray[19][42], dotarray[20][42], dotarray[21][42], dotarray[22][42], dotarray[23][42], dotarray[24][42], dotarray[25][42], dotarray[26][42], dotarray[27][42], dotarray[28][42], dotarray[29][42], dotarray[30][42], dotarray[31][42], dotarray[32][42], dotarray[33][42], dotarray[34][42], dotarray[35][42], dotarray[36][42], dotarray[37][42], dotarray[38][42], dotarray[39][42], dotarray[40][42], dotarray[41][42], dotarray[42][42], dotarray[43][42], dotarray[44][42], dotarray[45][42], dotarray[46][42], dotarray[47][42], dotarray[48][42], dotarray[49][42], dotarray[50][42], dotarray[51][42], dotarray[52][42], dotarray[53][42], dotarray[54][42], dotarray[55][42], dotarray[56][42], dotarray[57][42], dotarray[58][42], dotarray[59][42], dotarray[60][42], dotarray[61][42], dotarray[62][42], dotarray[63][42], dotarray[64][42], dotarray[65][42], dotarray[66][42], dotarray[67][42], dotarray[68][42], dotarray[69][42], dotarray[70][42], dotarray[71][42], dotarray[72][42], dotarray[73][42], dotarray[74][42], dotarray[75][42], dotarray[76][42], dotarray[77][42], dotarray[78][42], dotarray[79][42], dotarray[80][42], dotarray[81][42], dotarray[82][42], dotarray[83][42], dotarray[84][42], dotarray[85][42], dotarray[86][42], dotarray[87][42], dotarray[88][42], dotarray[89][42], dotarray[90][42], dotarray[91][42], dotarray[92][42], dotarray[93][42], dotarray[94][42], dotarray[95][42], dotarray[96][42], dotarray[97][42], dotarray[98][42], dotarray[99][42], dotarray[100][42], dotarray[101][42], dotarray[102][42], dotarray[103][42], dotarray[104][42], dotarray[105][42], dotarray[106][42], dotarray[107][42], dotarray[108][42], dotarray[109][42], dotarray[110][42], dotarray[111][42], dotarray[112][42], dotarray[113][42], dotarray[114][42], dotarray[115][42], dotarray[116][42], dotarray[117][42], dotarray[118][42], dotarray[119][42], dotarray[120][42], dotarray[121][42], dotarray[122][42], dotarray[123][42], dotarray[124][42], dotarray[125][42], dotarray[126][42], dotarray[127][42]};
assign dot_col_43 = {dotarray[0][43], dotarray[1][43], dotarray[2][43], dotarray[3][43], dotarray[4][43], dotarray[5][43], dotarray[6][43], dotarray[7][43], dotarray[8][43], dotarray[9][43], dotarray[10][43], dotarray[11][43], dotarray[12][43], dotarray[13][43], dotarray[14][43], dotarray[15][43], dotarray[16][43], dotarray[17][43], dotarray[18][43], dotarray[19][43], dotarray[20][43], dotarray[21][43], dotarray[22][43], dotarray[23][43], dotarray[24][43], dotarray[25][43], dotarray[26][43], dotarray[27][43], dotarray[28][43], dotarray[29][43], dotarray[30][43], dotarray[31][43], dotarray[32][43], dotarray[33][43], dotarray[34][43], dotarray[35][43], dotarray[36][43], dotarray[37][43], dotarray[38][43], dotarray[39][43], dotarray[40][43], dotarray[41][43], dotarray[42][43], dotarray[43][43], dotarray[44][43], dotarray[45][43], dotarray[46][43], dotarray[47][43], dotarray[48][43], dotarray[49][43], dotarray[50][43], dotarray[51][43], dotarray[52][43], dotarray[53][43], dotarray[54][43], dotarray[55][43], dotarray[56][43], dotarray[57][43], dotarray[58][43], dotarray[59][43], dotarray[60][43], dotarray[61][43], dotarray[62][43], dotarray[63][43], dotarray[64][43], dotarray[65][43], dotarray[66][43], dotarray[67][43], dotarray[68][43], dotarray[69][43], dotarray[70][43], dotarray[71][43], dotarray[72][43], dotarray[73][43], dotarray[74][43], dotarray[75][43], dotarray[76][43], dotarray[77][43], dotarray[78][43], dotarray[79][43], dotarray[80][43], dotarray[81][43], dotarray[82][43], dotarray[83][43], dotarray[84][43], dotarray[85][43], dotarray[86][43], dotarray[87][43], dotarray[88][43], dotarray[89][43], dotarray[90][43], dotarray[91][43], dotarray[92][43], dotarray[93][43], dotarray[94][43], dotarray[95][43], dotarray[96][43], dotarray[97][43], dotarray[98][43], dotarray[99][43], dotarray[100][43], dotarray[101][43], dotarray[102][43], dotarray[103][43], dotarray[104][43], dotarray[105][43], dotarray[106][43], dotarray[107][43], dotarray[108][43], dotarray[109][43], dotarray[110][43], dotarray[111][43], dotarray[112][43], dotarray[113][43], dotarray[114][43], dotarray[115][43], dotarray[116][43], dotarray[117][43], dotarray[118][43], dotarray[119][43], dotarray[120][43], dotarray[121][43], dotarray[122][43], dotarray[123][43], dotarray[124][43], dotarray[125][43], dotarray[126][43], dotarray[127][43]};
assign dot_col_44 = {dotarray[0][44], dotarray[1][44], dotarray[2][44], dotarray[3][44], dotarray[4][44], dotarray[5][44], dotarray[6][44], dotarray[7][44], dotarray[8][44], dotarray[9][44], dotarray[10][44], dotarray[11][44], dotarray[12][44], dotarray[13][44], dotarray[14][44], dotarray[15][44], dotarray[16][44], dotarray[17][44], dotarray[18][44], dotarray[19][44], dotarray[20][44], dotarray[21][44], dotarray[22][44], dotarray[23][44], dotarray[24][44], dotarray[25][44], dotarray[26][44], dotarray[27][44], dotarray[28][44], dotarray[29][44], dotarray[30][44], dotarray[31][44], dotarray[32][44], dotarray[33][44], dotarray[34][44], dotarray[35][44], dotarray[36][44], dotarray[37][44], dotarray[38][44], dotarray[39][44], dotarray[40][44], dotarray[41][44], dotarray[42][44], dotarray[43][44], dotarray[44][44], dotarray[45][44], dotarray[46][44], dotarray[47][44], dotarray[48][44], dotarray[49][44], dotarray[50][44], dotarray[51][44], dotarray[52][44], dotarray[53][44], dotarray[54][44], dotarray[55][44], dotarray[56][44], dotarray[57][44], dotarray[58][44], dotarray[59][44], dotarray[60][44], dotarray[61][44], dotarray[62][44], dotarray[63][44], dotarray[64][44], dotarray[65][44], dotarray[66][44], dotarray[67][44], dotarray[68][44], dotarray[69][44], dotarray[70][44], dotarray[71][44], dotarray[72][44], dotarray[73][44], dotarray[74][44], dotarray[75][44], dotarray[76][44], dotarray[77][44], dotarray[78][44], dotarray[79][44], dotarray[80][44], dotarray[81][44], dotarray[82][44], dotarray[83][44], dotarray[84][44], dotarray[85][44], dotarray[86][44], dotarray[87][44], dotarray[88][44], dotarray[89][44], dotarray[90][44], dotarray[91][44], dotarray[92][44], dotarray[93][44], dotarray[94][44], dotarray[95][44], dotarray[96][44], dotarray[97][44], dotarray[98][44], dotarray[99][44], dotarray[100][44], dotarray[101][44], dotarray[102][44], dotarray[103][44], dotarray[104][44], dotarray[105][44], dotarray[106][44], dotarray[107][44], dotarray[108][44], dotarray[109][44], dotarray[110][44], dotarray[111][44], dotarray[112][44], dotarray[113][44], dotarray[114][44], dotarray[115][44], dotarray[116][44], dotarray[117][44], dotarray[118][44], dotarray[119][44], dotarray[120][44], dotarray[121][44], dotarray[122][44], dotarray[123][44], dotarray[124][44], dotarray[125][44], dotarray[126][44], dotarray[127][44]};
assign dot_col_45 = {dotarray[0][45], dotarray[1][45], dotarray[2][45], dotarray[3][45], dotarray[4][45], dotarray[5][45], dotarray[6][45], dotarray[7][45], dotarray[8][45], dotarray[9][45], dotarray[10][45], dotarray[11][45], dotarray[12][45], dotarray[13][45], dotarray[14][45], dotarray[15][45], dotarray[16][45], dotarray[17][45], dotarray[18][45], dotarray[19][45], dotarray[20][45], dotarray[21][45], dotarray[22][45], dotarray[23][45], dotarray[24][45], dotarray[25][45], dotarray[26][45], dotarray[27][45], dotarray[28][45], dotarray[29][45], dotarray[30][45], dotarray[31][45], dotarray[32][45], dotarray[33][45], dotarray[34][45], dotarray[35][45], dotarray[36][45], dotarray[37][45], dotarray[38][45], dotarray[39][45], dotarray[40][45], dotarray[41][45], dotarray[42][45], dotarray[43][45], dotarray[44][45], dotarray[45][45], dotarray[46][45], dotarray[47][45], dotarray[48][45], dotarray[49][45], dotarray[50][45], dotarray[51][45], dotarray[52][45], dotarray[53][45], dotarray[54][45], dotarray[55][45], dotarray[56][45], dotarray[57][45], dotarray[58][45], dotarray[59][45], dotarray[60][45], dotarray[61][45], dotarray[62][45], dotarray[63][45], dotarray[64][45], dotarray[65][45], dotarray[66][45], dotarray[67][45], dotarray[68][45], dotarray[69][45], dotarray[70][45], dotarray[71][45], dotarray[72][45], dotarray[73][45], dotarray[74][45], dotarray[75][45], dotarray[76][45], dotarray[77][45], dotarray[78][45], dotarray[79][45], dotarray[80][45], dotarray[81][45], dotarray[82][45], dotarray[83][45], dotarray[84][45], dotarray[85][45], dotarray[86][45], dotarray[87][45], dotarray[88][45], dotarray[89][45], dotarray[90][45], dotarray[91][45], dotarray[92][45], dotarray[93][45], dotarray[94][45], dotarray[95][45], dotarray[96][45], dotarray[97][45], dotarray[98][45], dotarray[99][45], dotarray[100][45], dotarray[101][45], dotarray[102][45], dotarray[103][45], dotarray[104][45], dotarray[105][45], dotarray[106][45], dotarray[107][45], dotarray[108][45], dotarray[109][45], dotarray[110][45], dotarray[111][45], dotarray[112][45], dotarray[113][45], dotarray[114][45], dotarray[115][45], dotarray[116][45], dotarray[117][45], dotarray[118][45], dotarray[119][45], dotarray[120][45], dotarray[121][45], dotarray[122][45], dotarray[123][45], dotarray[124][45], dotarray[125][45], dotarray[126][45], dotarray[127][45]};
assign dot_col_46 = {dotarray[0][46], dotarray[1][46], dotarray[2][46], dotarray[3][46], dotarray[4][46], dotarray[5][46], dotarray[6][46], dotarray[7][46], dotarray[8][46], dotarray[9][46], dotarray[10][46], dotarray[11][46], dotarray[12][46], dotarray[13][46], dotarray[14][46], dotarray[15][46], dotarray[16][46], dotarray[17][46], dotarray[18][46], dotarray[19][46], dotarray[20][46], dotarray[21][46], dotarray[22][46], dotarray[23][46], dotarray[24][46], dotarray[25][46], dotarray[26][46], dotarray[27][46], dotarray[28][46], dotarray[29][46], dotarray[30][46], dotarray[31][46], dotarray[32][46], dotarray[33][46], dotarray[34][46], dotarray[35][46], dotarray[36][46], dotarray[37][46], dotarray[38][46], dotarray[39][46], dotarray[40][46], dotarray[41][46], dotarray[42][46], dotarray[43][46], dotarray[44][46], dotarray[45][46], dotarray[46][46], dotarray[47][46], dotarray[48][46], dotarray[49][46], dotarray[50][46], dotarray[51][46], dotarray[52][46], dotarray[53][46], dotarray[54][46], dotarray[55][46], dotarray[56][46], dotarray[57][46], dotarray[58][46], dotarray[59][46], dotarray[60][46], dotarray[61][46], dotarray[62][46], dotarray[63][46], dotarray[64][46], dotarray[65][46], dotarray[66][46], dotarray[67][46], dotarray[68][46], dotarray[69][46], dotarray[70][46], dotarray[71][46], dotarray[72][46], dotarray[73][46], dotarray[74][46], dotarray[75][46], dotarray[76][46], dotarray[77][46], dotarray[78][46], dotarray[79][46], dotarray[80][46], dotarray[81][46], dotarray[82][46], dotarray[83][46], dotarray[84][46], dotarray[85][46], dotarray[86][46], dotarray[87][46], dotarray[88][46], dotarray[89][46], dotarray[90][46], dotarray[91][46], dotarray[92][46], dotarray[93][46], dotarray[94][46], dotarray[95][46], dotarray[96][46], dotarray[97][46], dotarray[98][46], dotarray[99][46], dotarray[100][46], dotarray[101][46], dotarray[102][46], dotarray[103][46], dotarray[104][46], dotarray[105][46], dotarray[106][46], dotarray[107][46], dotarray[108][46], dotarray[109][46], dotarray[110][46], dotarray[111][46], dotarray[112][46], dotarray[113][46], dotarray[114][46], dotarray[115][46], dotarray[116][46], dotarray[117][46], dotarray[118][46], dotarray[119][46], dotarray[120][46], dotarray[121][46], dotarray[122][46], dotarray[123][46], dotarray[124][46], dotarray[125][46], dotarray[126][46], dotarray[127][46]};
assign dot_col_47 = {dotarray[0][47], dotarray[1][47], dotarray[2][47], dotarray[3][47], dotarray[4][47], dotarray[5][47], dotarray[6][47], dotarray[7][47], dotarray[8][47], dotarray[9][47], dotarray[10][47], dotarray[11][47], dotarray[12][47], dotarray[13][47], dotarray[14][47], dotarray[15][47], dotarray[16][47], dotarray[17][47], dotarray[18][47], dotarray[19][47], dotarray[20][47], dotarray[21][47], dotarray[22][47], dotarray[23][47], dotarray[24][47], dotarray[25][47], dotarray[26][47], dotarray[27][47], dotarray[28][47], dotarray[29][47], dotarray[30][47], dotarray[31][47], dotarray[32][47], dotarray[33][47], dotarray[34][47], dotarray[35][47], dotarray[36][47], dotarray[37][47], dotarray[38][47], dotarray[39][47], dotarray[40][47], dotarray[41][47], dotarray[42][47], dotarray[43][47], dotarray[44][47], dotarray[45][47], dotarray[46][47], dotarray[47][47], dotarray[48][47], dotarray[49][47], dotarray[50][47], dotarray[51][47], dotarray[52][47], dotarray[53][47], dotarray[54][47], dotarray[55][47], dotarray[56][47], dotarray[57][47], dotarray[58][47], dotarray[59][47], dotarray[60][47], dotarray[61][47], dotarray[62][47], dotarray[63][47], dotarray[64][47], dotarray[65][47], dotarray[66][47], dotarray[67][47], dotarray[68][47], dotarray[69][47], dotarray[70][47], dotarray[71][47], dotarray[72][47], dotarray[73][47], dotarray[74][47], dotarray[75][47], dotarray[76][47], dotarray[77][47], dotarray[78][47], dotarray[79][47], dotarray[80][47], dotarray[81][47], dotarray[82][47], dotarray[83][47], dotarray[84][47], dotarray[85][47], dotarray[86][47], dotarray[87][47], dotarray[88][47], dotarray[89][47], dotarray[90][47], dotarray[91][47], dotarray[92][47], dotarray[93][47], dotarray[94][47], dotarray[95][47], dotarray[96][47], dotarray[97][47], dotarray[98][47], dotarray[99][47], dotarray[100][47], dotarray[101][47], dotarray[102][47], dotarray[103][47], dotarray[104][47], dotarray[105][47], dotarray[106][47], dotarray[107][47], dotarray[108][47], dotarray[109][47], dotarray[110][47], dotarray[111][47], dotarray[112][47], dotarray[113][47], dotarray[114][47], dotarray[115][47], dotarray[116][47], dotarray[117][47], dotarray[118][47], dotarray[119][47], dotarray[120][47], dotarray[121][47], dotarray[122][47], dotarray[123][47], dotarray[124][47], dotarray[125][47], dotarray[126][47], dotarray[127][47]};
assign dot_col_48 = {dotarray[0][48], dotarray[1][48], dotarray[2][48], dotarray[3][48], dotarray[4][48], dotarray[5][48], dotarray[6][48], dotarray[7][48], dotarray[8][48], dotarray[9][48], dotarray[10][48], dotarray[11][48], dotarray[12][48], dotarray[13][48], dotarray[14][48], dotarray[15][48], dotarray[16][48], dotarray[17][48], dotarray[18][48], dotarray[19][48], dotarray[20][48], dotarray[21][48], dotarray[22][48], dotarray[23][48], dotarray[24][48], dotarray[25][48], dotarray[26][48], dotarray[27][48], dotarray[28][48], dotarray[29][48], dotarray[30][48], dotarray[31][48], dotarray[32][48], dotarray[33][48], dotarray[34][48], dotarray[35][48], dotarray[36][48], dotarray[37][48], dotarray[38][48], dotarray[39][48], dotarray[40][48], dotarray[41][48], dotarray[42][48], dotarray[43][48], dotarray[44][48], dotarray[45][48], dotarray[46][48], dotarray[47][48], dotarray[48][48], dotarray[49][48], dotarray[50][48], dotarray[51][48], dotarray[52][48], dotarray[53][48], dotarray[54][48], dotarray[55][48], dotarray[56][48], dotarray[57][48], dotarray[58][48], dotarray[59][48], dotarray[60][48], dotarray[61][48], dotarray[62][48], dotarray[63][48], dotarray[64][48], dotarray[65][48], dotarray[66][48], dotarray[67][48], dotarray[68][48], dotarray[69][48], dotarray[70][48], dotarray[71][48], dotarray[72][48], dotarray[73][48], dotarray[74][48], dotarray[75][48], dotarray[76][48], dotarray[77][48], dotarray[78][48], dotarray[79][48], dotarray[80][48], dotarray[81][48], dotarray[82][48], dotarray[83][48], dotarray[84][48], dotarray[85][48], dotarray[86][48], dotarray[87][48], dotarray[88][48], dotarray[89][48], dotarray[90][48], dotarray[91][48], dotarray[92][48], dotarray[93][48], dotarray[94][48], dotarray[95][48], dotarray[96][48], dotarray[97][48], dotarray[98][48], dotarray[99][48], dotarray[100][48], dotarray[101][48], dotarray[102][48], dotarray[103][48], dotarray[104][48], dotarray[105][48], dotarray[106][48], dotarray[107][48], dotarray[108][48], dotarray[109][48], dotarray[110][48], dotarray[111][48], dotarray[112][48], dotarray[113][48], dotarray[114][48], dotarray[115][48], dotarray[116][48], dotarray[117][48], dotarray[118][48], dotarray[119][48], dotarray[120][48], dotarray[121][48], dotarray[122][48], dotarray[123][48], dotarray[124][48], dotarray[125][48], dotarray[126][48], dotarray[127][48]};
assign dot_col_49 = {dotarray[0][49], dotarray[1][49], dotarray[2][49], dotarray[3][49], dotarray[4][49], dotarray[5][49], dotarray[6][49], dotarray[7][49], dotarray[8][49], dotarray[9][49], dotarray[10][49], dotarray[11][49], dotarray[12][49], dotarray[13][49], dotarray[14][49], dotarray[15][49], dotarray[16][49], dotarray[17][49], dotarray[18][49], dotarray[19][49], dotarray[20][49], dotarray[21][49], dotarray[22][49], dotarray[23][49], dotarray[24][49], dotarray[25][49], dotarray[26][49], dotarray[27][49], dotarray[28][49], dotarray[29][49], dotarray[30][49], dotarray[31][49], dotarray[32][49], dotarray[33][49], dotarray[34][49], dotarray[35][49], dotarray[36][49], dotarray[37][49], dotarray[38][49], dotarray[39][49], dotarray[40][49], dotarray[41][49], dotarray[42][49], dotarray[43][49], dotarray[44][49], dotarray[45][49], dotarray[46][49], dotarray[47][49], dotarray[48][49], dotarray[49][49], dotarray[50][49], dotarray[51][49], dotarray[52][49], dotarray[53][49], dotarray[54][49], dotarray[55][49], dotarray[56][49], dotarray[57][49], dotarray[58][49], dotarray[59][49], dotarray[60][49], dotarray[61][49], dotarray[62][49], dotarray[63][49], dotarray[64][49], dotarray[65][49], dotarray[66][49], dotarray[67][49], dotarray[68][49], dotarray[69][49], dotarray[70][49], dotarray[71][49], dotarray[72][49], dotarray[73][49], dotarray[74][49], dotarray[75][49], dotarray[76][49], dotarray[77][49], dotarray[78][49], dotarray[79][49], dotarray[80][49], dotarray[81][49], dotarray[82][49], dotarray[83][49], dotarray[84][49], dotarray[85][49], dotarray[86][49], dotarray[87][49], dotarray[88][49], dotarray[89][49], dotarray[90][49], dotarray[91][49], dotarray[92][49], dotarray[93][49], dotarray[94][49], dotarray[95][49], dotarray[96][49], dotarray[97][49], dotarray[98][49], dotarray[99][49], dotarray[100][49], dotarray[101][49], dotarray[102][49], dotarray[103][49], dotarray[104][49], dotarray[105][49], dotarray[106][49], dotarray[107][49], dotarray[108][49], dotarray[109][49], dotarray[110][49], dotarray[111][49], dotarray[112][49], dotarray[113][49], dotarray[114][49], dotarray[115][49], dotarray[116][49], dotarray[117][49], dotarray[118][49], dotarray[119][49], dotarray[120][49], dotarray[121][49], dotarray[122][49], dotarray[123][49], dotarray[124][49], dotarray[125][49], dotarray[126][49], dotarray[127][49]};
assign dot_col_50 = {dotarray[0][50], dotarray[1][50], dotarray[2][50], dotarray[3][50], dotarray[4][50], dotarray[5][50], dotarray[6][50], dotarray[7][50], dotarray[8][50], dotarray[9][50], dotarray[10][50], dotarray[11][50], dotarray[12][50], dotarray[13][50], dotarray[14][50], dotarray[15][50], dotarray[16][50], dotarray[17][50], dotarray[18][50], dotarray[19][50], dotarray[20][50], dotarray[21][50], dotarray[22][50], dotarray[23][50], dotarray[24][50], dotarray[25][50], dotarray[26][50], dotarray[27][50], dotarray[28][50], dotarray[29][50], dotarray[30][50], dotarray[31][50], dotarray[32][50], dotarray[33][50], dotarray[34][50], dotarray[35][50], dotarray[36][50], dotarray[37][50], dotarray[38][50], dotarray[39][50], dotarray[40][50], dotarray[41][50], dotarray[42][50], dotarray[43][50], dotarray[44][50], dotarray[45][50], dotarray[46][50], dotarray[47][50], dotarray[48][50], dotarray[49][50], dotarray[50][50], dotarray[51][50], dotarray[52][50], dotarray[53][50], dotarray[54][50], dotarray[55][50], dotarray[56][50], dotarray[57][50], dotarray[58][50], dotarray[59][50], dotarray[60][50], dotarray[61][50], dotarray[62][50], dotarray[63][50], dotarray[64][50], dotarray[65][50], dotarray[66][50], dotarray[67][50], dotarray[68][50], dotarray[69][50], dotarray[70][50], dotarray[71][50], dotarray[72][50], dotarray[73][50], dotarray[74][50], dotarray[75][50], dotarray[76][50], dotarray[77][50], dotarray[78][50], dotarray[79][50], dotarray[80][50], dotarray[81][50], dotarray[82][50], dotarray[83][50], dotarray[84][50], dotarray[85][50], dotarray[86][50], dotarray[87][50], dotarray[88][50], dotarray[89][50], dotarray[90][50], dotarray[91][50], dotarray[92][50], dotarray[93][50], dotarray[94][50], dotarray[95][50], dotarray[96][50], dotarray[97][50], dotarray[98][50], dotarray[99][50], dotarray[100][50], dotarray[101][50], dotarray[102][50], dotarray[103][50], dotarray[104][50], dotarray[105][50], dotarray[106][50], dotarray[107][50], dotarray[108][50], dotarray[109][50], dotarray[110][50], dotarray[111][50], dotarray[112][50], dotarray[113][50], dotarray[114][50], dotarray[115][50], dotarray[116][50], dotarray[117][50], dotarray[118][50], dotarray[119][50], dotarray[120][50], dotarray[121][50], dotarray[122][50], dotarray[123][50], dotarray[124][50], dotarray[125][50], dotarray[126][50], dotarray[127][50]};
assign dot_col_51 = {dotarray[0][51], dotarray[1][51], dotarray[2][51], dotarray[3][51], dotarray[4][51], dotarray[5][51], dotarray[6][51], dotarray[7][51], dotarray[8][51], dotarray[9][51], dotarray[10][51], dotarray[11][51], dotarray[12][51], dotarray[13][51], dotarray[14][51], dotarray[15][51], dotarray[16][51], dotarray[17][51], dotarray[18][51], dotarray[19][51], dotarray[20][51], dotarray[21][51], dotarray[22][51], dotarray[23][51], dotarray[24][51], dotarray[25][51], dotarray[26][51], dotarray[27][51], dotarray[28][51], dotarray[29][51], dotarray[30][51], dotarray[31][51], dotarray[32][51], dotarray[33][51], dotarray[34][51], dotarray[35][51], dotarray[36][51], dotarray[37][51], dotarray[38][51], dotarray[39][51], dotarray[40][51], dotarray[41][51], dotarray[42][51], dotarray[43][51], dotarray[44][51], dotarray[45][51], dotarray[46][51], dotarray[47][51], dotarray[48][51], dotarray[49][51], dotarray[50][51], dotarray[51][51], dotarray[52][51], dotarray[53][51], dotarray[54][51], dotarray[55][51], dotarray[56][51], dotarray[57][51], dotarray[58][51], dotarray[59][51], dotarray[60][51], dotarray[61][51], dotarray[62][51], dotarray[63][51], dotarray[64][51], dotarray[65][51], dotarray[66][51], dotarray[67][51], dotarray[68][51], dotarray[69][51], dotarray[70][51], dotarray[71][51], dotarray[72][51], dotarray[73][51], dotarray[74][51], dotarray[75][51], dotarray[76][51], dotarray[77][51], dotarray[78][51], dotarray[79][51], dotarray[80][51], dotarray[81][51], dotarray[82][51], dotarray[83][51], dotarray[84][51], dotarray[85][51], dotarray[86][51], dotarray[87][51], dotarray[88][51], dotarray[89][51], dotarray[90][51], dotarray[91][51], dotarray[92][51], dotarray[93][51], dotarray[94][51], dotarray[95][51], dotarray[96][51], dotarray[97][51], dotarray[98][51], dotarray[99][51], dotarray[100][51], dotarray[101][51], dotarray[102][51], dotarray[103][51], dotarray[104][51], dotarray[105][51], dotarray[106][51], dotarray[107][51], dotarray[108][51], dotarray[109][51], dotarray[110][51], dotarray[111][51], dotarray[112][51], dotarray[113][51], dotarray[114][51], dotarray[115][51], dotarray[116][51], dotarray[117][51], dotarray[118][51], dotarray[119][51], dotarray[120][51], dotarray[121][51], dotarray[122][51], dotarray[123][51], dotarray[124][51], dotarray[125][51], dotarray[126][51], dotarray[127][51]};
assign dot_col_52 = {dotarray[0][52], dotarray[1][52], dotarray[2][52], dotarray[3][52], dotarray[4][52], dotarray[5][52], dotarray[6][52], dotarray[7][52], dotarray[8][52], dotarray[9][52], dotarray[10][52], dotarray[11][52], dotarray[12][52], dotarray[13][52], dotarray[14][52], dotarray[15][52], dotarray[16][52], dotarray[17][52], dotarray[18][52], dotarray[19][52], dotarray[20][52], dotarray[21][52], dotarray[22][52], dotarray[23][52], dotarray[24][52], dotarray[25][52], dotarray[26][52], dotarray[27][52], dotarray[28][52], dotarray[29][52], dotarray[30][52], dotarray[31][52], dotarray[32][52], dotarray[33][52], dotarray[34][52], dotarray[35][52], dotarray[36][52], dotarray[37][52], dotarray[38][52], dotarray[39][52], dotarray[40][52], dotarray[41][52], dotarray[42][52], dotarray[43][52], dotarray[44][52], dotarray[45][52], dotarray[46][52], dotarray[47][52], dotarray[48][52], dotarray[49][52], dotarray[50][52], dotarray[51][52], dotarray[52][52], dotarray[53][52], dotarray[54][52], dotarray[55][52], dotarray[56][52], dotarray[57][52], dotarray[58][52], dotarray[59][52], dotarray[60][52], dotarray[61][52], dotarray[62][52], dotarray[63][52], dotarray[64][52], dotarray[65][52], dotarray[66][52], dotarray[67][52], dotarray[68][52], dotarray[69][52], dotarray[70][52], dotarray[71][52], dotarray[72][52], dotarray[73][52], dotarray[74][52], dotarray[75][52], dotarray[76][52], dotarray[77][52], dotarray[78][52], dotarray[79][52], dotarray[80][52], dotarray[81][52], dotarray[82][52], dotarray[83][52], dotarray[84][52], dotarray[85][52], dotarray[86][52], dotarray[87][52], dotarray[88][52], dotarray[89][52], dotarray[90][52], dotarray[91][52], dotarray[92][52], dotarray[93][52], dotarray[94][52], dotarray[95][52], dotarray[96][52], dotarray[97][52], dotarray[98][52], dotarray[99][52], dotarray[100][52], dotarray[101][52], dotarray[102][52], dotarray[103][52], dotarray[104][52], dotarray[105][52], dotarray[106][52], dotarray[107][52], dotarray[108][52], dotarray[109][52], dotarray[110][52], dotarray[111][52], dotarray[112][52], dotarray[113][52], dotarray[114][52], dotarray[115][52], dotarray[116][52], dotarray[117][52], dotarray[118][52], dotarray[119][52], dotarray[120][52], dotarray[121][52], dotarray[122][52], dotarray[123][52], dotarray[124][52], dotarray[125][52], dotarray[126][52], dotarray[127][52]};
assign dot_col_53 = {dotarray[0][53], dotarray[1][53], dotarray[2][53], dotarray[3][53], dotarray[4][53], dotarray[5][53], dotarray[6][53], dotarray[7][53], dotarray[8][53], dotarray[9][53], dotarray[10][53], dotarray[11][53], dotarray[12][53], dotarray[13][53], dotarray[14][53], dotarray[15][53], dotarray[16][53], dotarray[17][53], dotarray[18][53], dotarray[19][53], dotarray[20][53], dotarray[21][53], dotarray[22][53], dotarray[23][53], dotarray[24][53], dotarray[25][53], dotarray[26][53], dotarray[27][53], dotarray[28][53], dotarray[29][53], dotarray[30][53], dotarray[31][53], dotarray[32][53], dotarray[33][53], dotarray[34][53], dotarray[35][53], dotarray[36][53], dotarray[37][53], dotarray[38][53], dotarray[39][53], dotarray[40][53], dotarray[41][53], dotarray[42][53], dotarray[43][53], dotarray[44][53], dotarray[45][53], dotarray[46][53], dotarray[47][53], dotarray[48][53], dotarray[49][53], dotarray[50][53], dotarray[51][53], dotarray[52][53], dotarray[53][53], dotarray[54][53], dotarray[55][53], dotarray[56][53], dotarray[57][53], dotarray[58][53], dotarray[59][53], dotarray[60][53], dotarray[61][53], dotarray[62][53], dotarray[63][53], dotarray[64][53], dotarray[65][53], dotarray[66][53], dotarray[67][53], dotarray[68][53], dotarray[69][53], dotarray[70][53], dotarray[71][53], dotarray[72][53], dotarray[73][53], dotarray[74][53], dotarray[75][53], dotarray[76][53], dotarray[77][53], dotarray[78][53], dotarray[79][53], dotarray[80][53], dotarray[81][53], dotarray[82][53], dotarray[83][53], dotarray[84][53], dotarray[85][53], dotarray[86][53], dotarray[87][53], dotarray[88][53], dotarray[89][53], dotarray[90][53], dotarray[91][53], dotarray[92][53], dotarray[93][53], dotarray[94][53], dotarray[95][53], dotarray[96][53], dotarray[97][53], dotarray[98][53], dotarray[99][53], dotarray[100][53], dotarray[101][53], dotarray[102][53], dotarray[103][53], dotarray[104][53], dotarray[105][53], dotarray[106][53], dotarray[107][53], dotarray[108][53], dotarray[109][53], dotarray[110][53], dotarray[111][53], dotarray[112][53], dotarray[113][53], dotarray[114][53], dotarray[115][53], dotarray[116][53], dotarray[117][53], dotarray[118][53], dotarray[119][53], dotarray[120][53], dotarray[121][53], dotarray[122][53], dotarray[123][53], dotarray[124][53], dotarray[125][53], dotarray[126][53], dotarray[127][53]};
assign dot_col_54 = {dotarray[0][54], dotarray[1][54], dotarray[2][54], dotarray[3][54], dotarray[4][54], dotarray[5][54], dotarray[6][54], dotarray[7][54], dotarray[8][54], dotarray[9][54], dotarray[10][54], dotarray[11][54], dotarray[12][54], dotarray[13][54], dotarray[14][54], dotarray[15][54], dotarray[16][54], dotarray[17][54], dotarray[18][54], dotarray[19][54], dotarray[20][54], dotarray[21][54], dotarray[22][54], dotarray[23][54], dotarray[24][54], dotarray[25][54], dotarray[26][54], dotarray[27][54], dotarray[28][54], dotarray[29][54], dotarray[30][54], dotarray[31][54], dotarray[32][54], dotarray[33][54], dotarray[34][54], dotarray[35][54], dotarray[36][54], dotarray[37][54], dotarray[38][54], dotarray[39][54], dotarray[40][54], dotarray[41][54], dotarray[42][54], dotarray[43][54], dotarray[44][54], dotarray[45][54], dotarray[46][54], dotarray[47][54], dotarray[48][54], dotarray[49][54], dotarray[50][54], dotarray[51][54], dotarray[52][54], dotarray[53][54], dotarray[54][54], dotarray[55][54], dotarray[56][54], dotarray[57][54], dotarray[58][54], dotarray[59][54], dotarray[60][54], dotarray[61][54], dotarray[62][54], dotarray[63][54], dotarray[64][54], dotarray[65][54], dotarray[66][54], dotarray[67][54], dotarray[68][54], dotarray[69][54], dotarray[70][54], dotarray[71][54], dotarray[72][54], dotarray[73][54], dotarray[74][54], dotarray[75][54], dotarray[76][54], dotarray[77][54], dotarray[78][54], dotarray[79][54], dotarray[80][54], dotarray[81][54], dotarray[82][54], dotarray[83][54], dotarray[84][54], dotarray[85][54], dotarray[86][54], dotarray[87][54], dotarray[88][54], dotarray[89][54], dotarray[90][54], dotarray[91][54], dotarray[92][54], dotarray[93][54], dotarray[94][54], dotarray[95][54], dotarray[96][54], dotarray[97][54], dotarray[98][54], dotarray[99][54], dotarray[100][54], dotarray[101][54], dotarray[102][54], dotarray[103][54], dotarray[104][54], dotarray[105][54], dotarray[106][54], dotarray[107][54], dotarray[108][54], dotarray[109][54], dotarray[110][54], dotarray[111][54], dotarray[112][54], dotarray[113][54], dotarray[114][54], dotarray[115][54], dotarray[116][54], dotarray[117][54], dotarray[118][54], dotarray[119][54], dotarray[120][54], dotarray[121][54], dotarray[122][54], dotarray[123][54], dotarray[124][54], dotarray[125][54], dotarray[126][54], dotarray[127][54]};
assign dot_col_55 = {dotarray[0][55], dotarray[1][55], dotarray[2][55], dotarray[3][55], dotarray[4][55], dotarray[5][55], dotarray[6][55], dotarray[7][55], dotarray[8][55], dotarray[9][55], dotarray[10][55], dotarray[11][55], dotarray[12][55], dotarray[13][55], dotarray[14][55], dotarray[15][55], dotarray[16][55], dotarray[17][55], dotarray[18][55], dotarray[19][55], dotarray[20][55], dotarray[21][55], dotarray[22][55], dotarray[23][55], dotarray[24][55], dotarray[25][55], dotarray[26][55], dotarray[27][55], dotarray[28][55], dotarray[29][55], dotarray[30][55], dotarray[31][55], dotarray[32][55], dotarray[33][55], dotarray[34][55], dotarray[35][55], dotarray[36][55], dotarray[37][55], dotarray[38][55], dotarray[39][55], dotarray[40][55], dotarray[41][55], dotarray[42][55], dotarray[43][55], dotarray[44][55], dotarray[45][55], dotarray[46][55], dotarray[47][55], dotarray[48][55], dotarray[49][55], dotarray[50][55], dotarray[51][55], dotarray[52][55], dotarray[53][55], dotarray[54][55], dotarray[55][55], dotarray[56][55], dotarray[57][55], dotarray[58][55], dotarray[59][55], dotarray[60][55], dotarray[61][55], dotarray[62][55], dotarray[63][55], dotarray[64][55], dotarray[65][55], dotarray[66][55], dotarray[67][55], dotarray[68][55], dotarray[69][55], dotarray[70][55], dotarray[71][55], dotarray[72][55], dotarray[73][55], dotarray[74][55], dotarray[75][55], dotarray[76][55], dotarray[77][55], dotarray[78][55], dotarray[79][55], dotarray[80][55], dotarray[81][55], dotarray[82][55], dotarray[83][55], dotarray[84][55], dotarray[85][55], dotarray[86][55], dotarray[87][55], dotarray[88][55], dotarray[89][55], dotarray[90][55], dotarray[91][55], dotarray[92][55], dotarray[93][55], dotarray[94][55], dotarray[95][55], dotarray[96][55], dotarray[97][55], dotarray[98][55], dotarray[99][55], dotarray[100][55], dotarray[101][55], dotarray[102][55], dotarray[103][55], dotarray[104][55], dotarray[105][55], dotarray[106][55], dotarray[107][55], dotarray[108][55], dotarray[109][55], dotarray[110][55], dotarray[111][55], dotarray[112][55], dotarray[113][55], dotarray[114][55], dotarray[115][55], dotarray[116][55], dotarray[117][55], dotarray[118][55], dotarray[119][55], dotarray[120][55], dotarray[121][55], dotarray[122][55], dotarray[123][55], dotarray[124][55], dotarray[125][55], dotarray[126][55], dotarray[127][55]};
assign dot_col_56 = {dotarray[0][56], dotarray[1][56], dotarray[2][56], dotarray[3][56], dotarray[4][56], dotarray[5][56], dotarray[6][56], dotarray[7][56], dotarray[8][56], dotarray[9][56], dotarray[10][56], dotarray[11][56], dotarray[12][56], dotarray[13][56], dotarray[14][56], dotarray[15][56], dotarray[16][56], dotarray[17][56], dotarray[18][56], dotarray[19][56], dotarray[20][56], dotarray[21][56], dotarray[22][56], dotarray[23][56], dotarray[24][56], dotarray[25][56], dotarray[26][56], dotarray[27][56], dotarray[28][56], dotarray[29][56], dotarray[30][56], dotarray[31][56], dotarray[32][56], dotarray[33][56], dotarray[34][56], dotarray[35][56], dotarray[36][56], dotarray[37][56], dotarray[38][56], dotarray[39][56], dotarray[40][56], dotarray[41][56], dotarray[42][56], dotarray[43][56], dotarray[44][56], dotarray[45][56], dotarray[46][56], dotarray[47][56], dotarray[48][56], dotarray[49][56], dotarray[50][56], dotarray[51][56], dotarray[52][56], dotarray[53][56], dotarray[54][56], dotarray[55][56], dotarray[56][56], dotarray[57][56], dotarray[58][56], dotarray[59][56], dotarray[60][56], dotarray[61][56], dotarray[62][56], dotarray[63][56], dotarray[64][56], dotarray[65][56], dotarray[66][56], dotarray[67][56], dotarray[68][56], dotarray[69][56], dotarray[70][56], dotarray[71][56], dotarray[72][56], dotarray[73][56], dotarray[74][56], dotarray[75][56], dotarray[76][56], dotarray[77][56], dotarray[78][56], dotarray[79][56], dotarray[80][56], dotarray[81][56], dotarray[82][56], dotarray[83][56], dotarray[84][56], dotarray[85][56], dotarray[86][56], dotarray[87][56], dotarray[88][56], dotarray[89][56], dotarray[90][56], dotarray[91][56], dotarray[92][56], dotarray[93][56], dotarray[94][56], dotarray[95][56], dotarray[96][56], dotarray[97][56], dotarray[98][56], dotarray[99][56], dotarray[100][56], dotarray[101][56], dotarray[102][56], dotarray[103][56], dotarray[104][56], dotarray[105][56], dotarray[106][56], dotarray[107][56], dotarray[108][56], dotarray[109][56], dotarray[110][56], dotarray[111][56], dotarray[112][56], dotarray[113][56], dotarray[114][56], dotarray[115][56], dotarray[116][56], dotarray[117][56], dotarray[118][56], dotarray[119][56], dotarray[120][56], dotarray[121][56], dotarray[122][56], dotarray[123][56], dotarray[124][56], dotarray[125][56], dotarray[126][56], dotarray[127][56]};
assign dot_col_57 = {dotarray[0][57], dotarray[1][57], dotarray[2][57], dotarray[3][57], dotarray[4][57], dotarray[5][57], dotarray[6][57], dotarray[7][57], dotarray[8][57], dotarray[9][57], dotarray[10][57], dotarray[11][57], dotarray[12][57], dotarray[13][57], dotarray[14][57], dotarray[15][57], dotarray[16][57], dotarray[17][57], dotarray[18][57], dotarray[19][57], dotarray[20][57], dotarray[21][57], dotarray[22][57], dotarray[23][57], dotarray[24][57], dotarray[25][57], dotarray[26][57], dotarray[27][57], dotarray[28][57], dotarray[29][57], dotarray[30][57], dotarray[31][57], dotarray[32][57], dotarray[33][57], dotarray[34][57], dotarray[35][57], dotarray[36][57], dotarray[37][57], dotarray[38][57], dotarray[39][57], dotarray[40][57], dotarray[41][57], dotarray[42][57], dotarray[43][57], dotarray[44][57], dotarray[45][57], dotarray[46][57], dotarray[47][57], dotarray[48][57], dotarray[49][57], dotarray[50][57], dotarray[51][57], dotarray[52][57], dotarray[53][57], dotarray[54][57], dotarray[55][57], dotarray[56][57], dotarray[57][57], dotarray[58][57], dotarray[59][57], dotarray[60][57], dotarray[61][57], dotarray[62][57], dotarray[63][57], dotarray[64][57], dotarray[65][57], dotarray[66][57], dotarray[67][57], dotarray[68][57], dotarray[69][57], dotarray[70][57], dotarray[71][57], dotarray[72][57], dotarray[73][57], dotarray[74][57], dotarray[75][57], dotarray[76][57], dotarray[77][57], dotarray[78][57], dotarray[79][57], dotarray[80][57], dotarray[81][57], dotarray[82][57], dotarray[83][57], dotarray[84][57], dotarray[85][57], dotarray[86][57], dotarray[87][57], dotarray[88][57], dotarray[89][57], dotarray[90][57], dotarray[91][57], dotarray[92][57], dotarray[93][57], dotarray[94][57], dotarray[95][57], dotarray[96][57], dotarray[97][57], dotarray[98][57], dotarray[99][57], dotarray[100][57], dotarray[101][57], dotarray[102][57], dotarray[103][57], dotarray[104][57], dotarray[105][57], dotarray[106][57], dotarray[107][57], dotarray[108][57], dotarray[109][57], dotarray[110][57], dotarray[111][57], dotarray[112][57], dotarray[113][57], dotarray[114][57], dotarray[115][57], dotarray[116][57], dotarray[117][57], dotarray[118][57], dotarray[119][57], dotarray[120][57], dotarray[121][57], dotarray[122][57], dotarray[123][57], dotarray[124][57], dotarray[125][57], dotarray[126][57], dotarray[127][57]};
assign dot_col_58 = {dotarray[0][58], dotarray[1][58], dotarray[2][58], dotarray[3][58], dotarray[4][58], dotarray[5][58], dotarray[6][58], dotarray[7][58], dotarray[8][58], dotarray[9][58], dotarray[10][58], dotarray[11][58], dotarray[12][58], dotarray[13][58], dotarray[14][58], dotarray[15][58], dotarray[16][58], dotarray[17][58], dotarray[18][58], dotarray[19][58], dotarray[20][58], dotarray[21][58], dotarray[22][58], dotarray[23][58], dotarray[24][58], dotarray[25][58], dotarray[26][58], dotarray[27][58], dotarray[28][58], dotarray[29][58], dotarray[30][58], dotarray[31][58], dotarray[32][58], dotarray[33][58], dotarray[34][58], dotarray[35][58], dotarray[36][58], dotarray[37][58], dotarray[38][58], dotarray[39][58], dotarray[40][58], dotarray[41][58], dotarray[42][58], dotarray[43][58], dotarray[44][58], dotarray[45][58], dotarray[46][58], dotarray[47][58], dotarray[48][58], dotarray[49][58], dotarray[50][58], dotarray[51][58], dotarray[52][58], dotarray[53][58], dotarray[54][58], dotarray[55][58], dotarray[56][58], dotarray[57][58], dotarray[58][58], dotarray[59][58], dotarray[60][58], dotarray[61][58], dotarray[62][58], dotarray[63][58], dotarray[64][58], dotarray[65][58], dotarray[66][58], dotarray[67][58], dotarray[68][58], dotarray[69][58], dotarray[70][58], dotarray[71][58], dotarray[72][58], dotarray[73][58], dotarray[74][58], dotarray[75][58], dotarray[76][58], dotarray[77][58], dotarray[78][58], dotarray[79][58], dotarray[80][58], dotarray[81][58], dotarray[82][58], dotarray[83][58], dotarray[84][58], dotarray[85][58], dotarray[86][58], dotarray[87][58], dotarray[88][58], dotarray[89][58], dotarray[90][58], dotarray[91][58], dotarray[92][58], dotarray[93][58], dotarray[94][58], dotarray[95][58], dotarray[96][58], dotarray[97][58], dotarray[98][58], dotarray[99][58], dotarray[100][58], dotarray[101][58], dotarray[102][58], dotarray[103][58], dotarray[104][58], dotarray[105][58], dotarray[106][58], dotarray[107][58], dotarray[108][58], dotarray[109][58], dotarray[110][58], dotarray[111][58], dotarray[112][58], dotarray[113][58], dotarray[114][58], dotarray[115][58], dotarray[116][58], dotarray[117][58], dotarray[118][58], dotarray[119][58], dotarray[120][58], dotarray[121][58], dotarray[122][58], dotarray[123][58], dotarray[124][58], dotarray[125][58], dotarray[126][58], dotarray[127][58]};
assign dot_col_59 = {dotarray[0][59], dotarray[1][59], dotarray[2][59], dotarray[3][59], dotarray[4][59], dotarray[5][59], dotarray[6][59], dotarray[7][59], dotarray[8][59], dotarray[9][59], dotarray[10][59], dotarray[11][59], dotarray[12][59], dotarray[13][59], dotarray[14][59], dotarray[15][59], dotarray[16][59], dotarray[17][59], dotarray[18][59], dotarray[19][59], dotarray[20][59], dotarray[21][59], dotarray[22][59], dotarray[23][59], dotarray[24][59], dotarray[25][59], dotarray[26][59], dotarray[27][59], dotarray[28][59], dotarray[29][59], dotarray[30][59], dotarray[31][59], dotarray[32][59], dotarray[33][59], dotarray[34][59], dotarray[35][59], dotarray[36][59], dotarray[37][59], dotarray[38][59], dotarray[39][59], dotarray[40][59], dotarray[41][59], dotarray[42][59], dotarray[43][59], dotarray[44][59], dotarray[45][59], dotarray[46][59], dotarray[47][59], dotarray[48][59], dotarray[49][59], dotarray[50][59], dotarray[51][59], dotarray[52][59], dotarray[53][59], dotarray[54][59], dotarray[55][59], dotarray[56][59], dotarray[57][59], dotarray[58][59], dotarray[59][59], dotarray[60][59], dotarray[61][59], dotarray[62][59], dotarray[63][59], dotarray[64][59], dotarray[65][59], dotarray[66][59], dotarray[67][59], dotarray[68][59], dotarray[69][59], dotarray[70][59], dotarray[71][59], dotarray[72][59], dotarray[73][59], dotarray[74][59], dotarray[75][59], dotarray[76][59], dotarray[77][59], dotarray[78][59], dotarray[79][59], dotarray[80][59], dotarray[81][59], dotarray[82][59], dotarray[83][59], dotarray[84][59], dotarray[85][59], dotarray[86][59], dotarray[87][59], dotarray[88][59], dotarray[89][59], dotarray[90][59], dotarray[91][59], dotarray[92][59], dotarray[93][59], dotarray[94][59], dotarray[95][59], dotarray[96][59], dotarray[97][59], dotarray[98][59], dotarray[99][59], dotarray[100][59], dotarray[101][59], dotarray[102][59], dotarray[103][59], dotarray[104][59], dotarray[105][59], dotarray[106][59], dotarray[107][59], dotarray[108][59], dotarray[109][59], dotarray[110][59], dotarray[111][59], dotarray[112][59], dotarray[113][59], dotarray[114][59], dotarray[115][59], dotarray[116][59], dotarray[117][59], dotarray[118][59], dotarray[119][59], dotarray[120][59], dotarray[121][59], dotarray[122][59], dotarray[123][59], dotarray[124][59], dotarray[125][59], dotarray[126][59], dotarray[127][59]};
assign dot_col_60 = {dotarray[0][60], dotarray[1][60], dotarray[2][60], dotarray[3][60], dotarray[4][60], dotarray[5][60], dotarray[6][60], dotarray[7][60], dotarray[8][60], dotarray[9][60], dotarray[10][60], dotarray[11][60], dotarray[12][60], dotarray[13][60], dotarray[14][60], dotarray[15][60], dotarray[16][60], dotarray[17][60], dotarray[18][60], dotarray[19][60], dotarray[20][60], dotarray[21][60], dotarray[22][60], dotarray[23][60], dotarray[24][60], dotarray[25][60], dotarray[26][60], dotarray[27][60], dotarray[28][60], dotarray[29][60], dotarray[30][60], dotarray[31][60], dotarray[32][60], dotarray[33][60], dotarray[34][60], dotarray[35][60], dotarray[36][60], dotarray[37][60], dotarray[38][60], dotarray[39][60], dotarray[40][60], dotarray[41][60], dotarray[42][60], dotarray[43][60], dotarray[44][60], dotarray[45][60], dotarray[46][60], dotarray[47][60], dotarray[48][60], dotarray[49][60], dotarray[50][60], dotarray[51][60], dotarray[52][60], dotarray[53][60], dotarray[54][60], dotarray[55][60], dotarray[56][60], dotarray[57][60], dotarray[58][60], dotarray[59][60], dotarray[60][60], dotarray[61][60], dotarray[62][60], dotarray[63][60], dotarray[64][60], dotarray[65][60], dotarray[66][60], dotarray[67][60], dotarray[68][60], dotarray[69][60], dotarray[70][60], dotarray[71][60], dotarray[72][60], dotarray[73][60], dotarray[74][60], dotarray[75][60], dotarray[76][60], dotarray[77][60], dotarray[78][60], dotarray[79][60], dotarray[80][60], dotarray[81][60], dotarray[82][60], dotarray[83][60], dotarray[84][60], dotarray[85][60], dotarray[86][60], dotarray[87][60], dotarray[88][60], dotarray[89][60], dotarray[90][60], dotarray[91][60], dotarray[92][60], dotarray[93][60], dotarray[94][60], dotarray[95][60], dotarray[96][60], dotarray[97][60], dotarray[98][60], dotarray[99][60], dotarray[100][60], dotarray[101][60], dotarray[102][60], dotarray[103][60], dotarray[104][60], dotarray[105][60], dotarray[106][60], dotarray[107][60], dotarray[108][60], dotarray[109][60], dotarray[110][60], dotarray[111][60], dotarray[112][60], dotarray[113][60], dotarray[114][60], dotarray[115][60], dotarray[116][60], dotarray[117][60], dotarray[118][60], dotarray[119][60], dotarray[120][60], dotarray[121][60], dotarray[122][60], dotarray[123][60], dotarray[124][60], dotarray[125][60], dotarray[126][60], dotarray[127][60]};
assign dot_col_61 = {dotarray[0][61], dotarray[1][61], dotarray[2][61], dotarray[3][61], dotarray[4][61], dotarray[5][61], dotarray[6][61], dotarray[7][61], dotarray[8][61], dotarray[9][61], dotarray[10][61], dotarray[11][61], dotarray[12][61], dotarray[13][61], dotarray[14][61], dotarray[15][61], dotarray[16][61], dotarray[17][61], dotarray[18][61], dotarray[19][61], dotarray[20][61], dotarray[21][61], dotarray[22][61], dotarray[23][61], dotarray[24][61], dotarray[25][61], dotarray[26][61], dotarray[27][61], dotarray[28][61], dotarray[29][61], dotarray[30][61], dotarray[31][61], dotarray[32][61], dotarray[33][61], dotarray[34][61], dotarray[35][61], dotarray[36][61], dotarray[37][61], dotarray[38][61], dotarray[39][61], dotarray[40][61], dotarray[41][61], dotarray[42][61], dotarray[43][61], dotarray[44][61], dotarray[45][61], dotarray[46][61], dotarray[47][61], dotarray[48][61], dotarray[49][61], dotarray[50][61], dotarray[51][61], dotarray[52][61], dotarray[53][61], dotarray[54][61], dotarray[55][61], dotarray[56][61], dotarray[57][61], dotarray[58][61], dotarray[59][61], dotarray[60][61], dotarray[61][61], dotarray[62][61], dotarray[63][61], dotarray[64][61], dotarray[65][61], dotarray[66][61], dotarray[67][61], dotarray[68][61], dotarray[69][61], dotarray[70][61], dotarray[71][61], dotarray[72][61], dotarray[73][61], dotarray[74][61], dotarray[75][61], dotarray[76][61], dotarray[77][61], dotarray[78][61], dotarray[79][61], dotarray[80][61], dotarray[81][61], dotarray[82][61], dotarray[83][61], dotarray[84][61], dotarray[85][61], dotarray[86][61], dotarray[87][61], dotarray[88][61], dotarray[89][61], dotarray[90][61], dotarray[91][61], dotarray[92][61], dotarray[93][61], dotarray[94][61], dotarray[95][61], dotarray[96][61], dotarray[97][61], dotarray[98][61], dotarray[99][61], dotarray[100][61], dotarray[101][61], dotarray[102][61], dotarray[103][61], dotarray[104][61], dotarray[105][61], dotarray[106][61], dotarray[107][61], dotarray[108][61], dotarray[109][61], dotarray[110][61], dotarray[111][61], dotarray[112][61], dotarray[113][61], dotarray[114][61], dotarray[115][61], dotarray[116][61], dotarray[117][61], dotarray[118][61], dotarray[119][61], dotarray[120][61], dotarray[121][61], dotarray[122][61], dotarray[123][61], dotarray[124][61], dotarray[125][61], dotarray[126][61], dotarray[127][61]};
assign dot_col_62 = {dotarray[0][62], dotarray[1][62], dotarray[2][62], dotarray[3][62], dotarray[4][62], dotarray[5][62], dotarray[6][62], dotarray[7][62], dotarray[8][62], dotarray[9][62], dotarray[10][62], dotarray[11][62], dotarray[12][62], dotarray[13][62], dotarray[14][62], dotarray[15][62], dotarray[16][62], dotarray[17][62], dotarray[18][62], dotarray[19][62], dotarray[20][62], dotarray[21][62], dotarray[22][62], dotarray[23][62], dotarray[24][62], dotarray[25][62], dotarray[26][62], dotarray[27][62], dotarray[28][62], dotarray[29][62], dotarray[30][62], dotarray[31][62], dotarray[32][62], dotarray[33][62], dotarray[34][62], dotarray[35][62], dotarray[36][62], dotarray[37][62], dotarray[38][62], dotarray[39][62], dotarray[40][62], dotarray[41][62], dotarray[42][62], dotarray[43][62], dotarray[44][62], dotarray[45][62], dotarray[46][62], dotarray[47][62], dotarray[48][62], dotarray[49][62], dotarray[50][62], dotarray[51][62], dotarray[52][62], dotarray[53][62], dotarray[54][62], dotarray[55][62], dotarray[56][62], dotarray[57][62], dotarray[58][62], dotarray[59][62], dotarray[60][62], dotarray[61][62], dotarray[62][62], dotarray[63][62], dotarray[64][62], dotarray[65][62], dotarray[66][62], dotarray[67][62], dotarray[68][62], dotarray[69][62], dotarray[70][62], dotarray[71][62], dotarray[72][62], dotarray[73][62], dotarray[74][62], dotarray[75][62], dotarray[76][62], dotarray[77][62], dotarray[78][62], dotarray[79][62], dotarray[80][62], dotarray[81][62], dotarray[82][62], dotarray[83][62], dotarray[84][62], dotarray[85][62], dotarray[86][62], dotarray[87][62], dotarray[88][62], dotarray[89][62], dotarray[90][62], dotarray[91][62], dotarray[92][62], dotarray[93][62], dotarray[94][62], dotarray[95][62], dotarray[96][62], dotarray[97][62], dotarray[98][62], dotarray[99][62], dotarray[100][62], dotarray[101][62], dotarray[102][62], dotarray[103][62], dotarray[104][62], dotarray[105][62], dotarray[106][62], dotarray[107][62], dotarray[108][62], dotarray[109][62], dotarray[110][62], dotarray[111][62], dotarray[112][62], dotarray[113][62], dotarray[114][62], dotarray[115][62], dotarray[116][62], dotarray[117][62], dotarray[118][62], dotarray[119][62], dotarray[120][62], dotarray[121][62], dotarray[122][62], dotarray[123][62], dotarray[124][62], dotarray[125][62], dotarray[126][62], dotarray[127][62]};
assign dot_col_63 = {dotarray[0][63], dotarray[1][63], dotarray[2][63], dotarray[3][63], dotarray[4][63], dotarray[5][63], dotarray[6][63], dotarray[7][63], dotarray[8][63], dotarray[9][63], dotarray[10][63], dotarray[11][63], dotarray[12][63], dotarray[13][63], dotarray[14][63], dotarray[15][63], dotarray[16][63], dotarray[17][63], dotarray[18][63], dotarray[19][63], dotarray[20][63], dotarray[21][63], dotarray[22][63], dotarray[23][63], dotarray[24][63], dotarray[25][63], dotarray[26][63], dotarray[27][63], dotarray[28][63], dotarray[29][63], dotarray[30][63], dotarray[31][63], dotarray[32][63], dotarray[33][63], dotarray[34][63], dotarray[35][63], dotarray[36][63], dotarray[37][63], dotarray[38][63], dotarray[39][63], dotarray[40][63], dotarray[41][63], dotarray[42][63], dotarray[43][63], dotarray[44][63], dotarray[45][63], dotarray[46][63], dotarray[47][63], dotarray[48][63], dotarray[49][63], dotarray[50][63], dotarray[51][63], dotarray[52][63], dotarray[53][63], dotarray[54][63], dotarray[55][63], dotarray[56][63], dotarray[57][63], dotarray[58][63], dotarray[59][63], dotarray[60][63], dotarray[61][63], dotarray[62][63], dotarray[63][63], dotarray[64][63], dotarray[65][63], dotarray[66][63], dotarray[67][63], dotarray[68][63], dotarray[69][63], dotarray[70][63], dotarray[71][63], dotarray[72][63], dotarray[73][63], dotarray[74][63], dotarray[75][63], dotarray[76][63], dotarray[77][63], dotarray[78][63], dotarray[79][63], dotarray[80][63], dotarray[81][63], dotarray[82][63], dotarray[83][63], dotarray[84][63], dotarray[85][63], dotarray[86][63], dotarray[87][63], dotarray[88][63], dotarray[89][63], dotarray[90][63], dotarray[91][63], dotarray[92][63], dotarray[93][63], dotarray[94][63], dotarray[95][63], dotarray[96][63], dotarray[97][63], dotarray[98][63], dotarray[99][63], dotarray[100][63], dotarray[101][63], dotarray[102][63], dotarray[103][63], dotarray[104][63], dotarray[105][63], dotarray[106][63], dotarray[107][63], dotarray[108][63], dotarray[109][63], dotarray[110][63], dotarray[111][63], dotarray[112][63], dotarray[113][63], dotarray[114][63], dotarray[115][63], dotarray[116][63], dotarray[117][63], dotarray[118][63], dotarray[119][63], dotarray[120][63], dotarray[121][63], dotarray[122][63], dotarray[123][63], dotarray[124][63], dotarray[125][63], dotarray[126][63], dotarray[127][63]};
assign dot_col_64 = {dotarray[0][64], dotarray[1][64], dotarray[2][64], dotarray[3][64], dotarray[4][64], dotarray[5][64], dotarray[6][64], dotarray[7][64], dotarray[8][64], dotarray[9][64], dotarray[10][64], dotarray[11][64], dotarray[12][64], dotarray[13][64], dotarray[14][64], dotarray[15][64], dotarray[16][64], dotarray[17][64], dotarray[18][64], dotarray[19][64], dotarray[20][64], dotarray[21][64], dotarray[22][64], dotarray[23][64], dotarray[24][64], dotarray[25][64], dotarray[26][64], dotarray[27][64], dotarray[28][64], dotarray[29][64], dotarray[30][64], dotarray[31][64], dotarray[32][64], dotarray[33][64], dotarray[34][64], dotarray[35][64], dotarray[36][64], dotarray[37][64], dotarray[38][64], dotarray[39][64], dotarray[40][64], dotarray[41][64], dotarray[42][64], dotarray[43][64], dotarray[44][64], dotarray[45][64], dotarray[46][64], dotarray[47][64], dotarray[48][64], dotarray[49][64], dotarray[50][64], dotarray[51][64], dotarray[52][64], dotarray[53][64], dotarray[54][64], dotarray[55][64], dotarray[56][64], dotarray[57][64], dotarray[58][64], dotarray[59][64], dotarray[60][64], dotarray[61][64], dotarray[62][64], dotarray[63][64], dotarray[64][64], dotarray[65][64], dotarray[66][64], dotarray[67][64], dotarray[68][64], dotarray[69][64], dotarray[70][64], dotarray[71][64], dotarray[72][64], dotarray[73][64], dotarray[74][64], dotarray[75][64], dotarray[76][64], dotarray[77][64], dotarray[78][64], dotarray[79][64], dotarray[80][64], dotarray[81][64], dotarray[82][64], dotarray[83][64], dotarray[84][64], dotarray[85][64], dotarray[86][64], dotarray[87][64], dotarray[88][64], dotarray[89][64], dotarray[90][64], dotarray[91][64], dotarray[92][64], dotarray[93][64], dotarray[94][64], dotarray[95][64], dotarray[96][64], dotarray[97][64], dotarray[98][64], dotarray[99][64], dotarray[100][64], dotarray[101][64], dotarray[102][64], dotarray[103][64], dotarray[104][64], dotarray[105][64], dotarray[106][64], dotarray[107][64], dotarray[108][64], dotarray[109][64], dotarray[110][64], dotarray[111][64], dotarray[112][64], dotarray[113][64], dotarray[114][64], dotarray[115][64], dotarray[116][64], dotarray[117][64], dotarray[118][64], dotarray[119][64], dotarray[120][64], dotarray[121][64], dotarray[122][64], dotarray[123][64], dotarray[124][64], dotarray[125][64], dotarray[126][64], dotarray[127][64]};
assign dot_col_65 = {dotarray[0][65], dotarray[1][65], dotarray[2][65], dotarray[3][65], dotarray[4][65], dotarray[5][65], dotarray[6][65], dotarray[7][65], dotarray[8][65], dotarray[9][65], dotarray[10][65], dotarray[11][65], dotarray[12][65], dotarray[13][65], dotarray[14][65], dotarray[15][65], dotarray[16][65], dotarray[17][65], dotarray[18][65], dotarray[19][65], dotarray[20][65], dotarray[21][65], dotarray[22][65], dotarray[23][65], dotarray[24][65], dotarray[25][65], dotarray[26][65], dotarray[27][65], dotarray[28][65], dotarray[29][65], dotarray[30][65], dotarray[31][65], dotarray[32][65], dotarray[33][65], dotarray[34][65], dotarray[35][65], dotarray[36][65], dotarray[37][65], dotarray[38][65], dotarray[39][65], dotarray[40][65], dotarray[41][65], dotarray[42][65], dotarray[43][65], dotarray[44][65], dotarray[45][65], dotarray[46][65], dotarray[47][65], dotarray[48][65], dotarray[49][65], dotarray[50][65], dotarray[51][65], dotarray[52][65], dotarray[53][65], dotarray[54][65], dotarray[55][65], dotarray[56][65], dotarray[57][65], dotarray[58][65], dotarray[59][65], dotarray[60][65], dotarray[61][65], dotarray[62][65], dotarray[63][65], dotarray[64][65], dotarray[65][65], dotarray[66][65], dotarray[67][65], dotarray[68][65], dotarray[69][65], dotarray[70][65], dotarray[71][65], dotarray[72][65], dotarray[73][65], dotarray[74][65], dotarray[75][65], dotarray[76][65], dotarray[77][65], dotarray[78][65], dotarray[79][65], dotarray[80][65], dotarray[81][65], dotarray[82][65], dotarray[83][65], dotarray[84][65], dotarray[85][65], dotarray[86][65], dotarray[87][65], dotarray[88][65], dotarray[89][65], dotarray[90][65], dotarray[91][65], dotarray[92][65], dotarray[93][65], dotarray[94][65], dotarray[95][65], dotarray[96][65], dotarray[97][65], dotarray[98][65], dotarray[99][65], dotarray[100][65], dotarray[101][65], dotarray[102][65], dotarray[103][65], dotarray[104][65], dotarray[105][65], dotarray[106][65], dotarray[107][65], dotarray[108][65], dotarray[109][65], dotarray[110][65], dotarray[111][65], dotarray[112][65], dotarray[113][65], dotarray[114][65], dotarray[115][65], dotarray[116][65], dotarray[117][65], dotarray[118][65], dotarray[119][65], dotarray[120][65], dotarray[121][65], dotarray[122][65], dotarray[123][65], dotarray[124][65], dotarray[125][65], dotarray[126][65], dotarray[127][65]};
assign dot_col_66 = {dotarray[0][66], dotarray[1][66], dotarray[2][66], dotarray[3][66], dotarray[4][66], dotarray[5][66], dotarray[6][66], dotarray[7][66], dotarray[8][66], dotarray[9][66], dotarray[10][66], dotarray[11][66], dotarray[12][66], dotarray[13][66], dotarray[14][66], dotarray[15][66], dotarray[16][66], dotarray[17][66], dotarray[18][66], dotarray[19][66], dotarray[20][66], dotarray[21][66], dotarray[22][66], dotarray[23][66], dotarray[24][66], dotarray[25][66], dotarray[26][66], dotarray[27][66], dotarray[28][66], dotarray[29][66], dotarray[30][66], dotarray[31][66], dotarray[32][66], dotarray[33][66], dotarray[34][66], dotarray[35][66], dotarray[36][66], dotarray[37][66], dotarray[38][66], dotarray[39][66], dotarray[40][66], dotarray[41][66], dotarray[42][66], dotarray[43][66], dotarray[44][66], dotarray[45][66], dotarray[46][66], dotarray[47][66], dotarray[48][66], dotarray[49][66], dotarray[50][66], dotarray[51][66], dotarray[52][66], dotarray[53][66], dotarray[54][66], dotarray[55][66], dotarray[56][66], dotarray[57][66], dotarray[58][66], dotarray[59][66], dotarray[60][66], dotarray[61][66], dotarray[62][66], dotarray[63][66], dotarray[64][66], dotarray[65][66], dotarray[66][66], dotarray[67][66], dotarray[68][66], dotarray[69][66], dotarray[70][66], dotarray[71][66], dotarray[72][66], dotarray[73][66], dotarray[74][66], dotarray[75][66], dotarray[76][66], dotarray[77][66], dotarray[78][66], dotarray[79][66], dotarray[80][66], dotarray[81][66], dotarray[82][66], dotarray[83][66], dotarray[84][66], dotarray[85][66], dotarray[86][66], dotarray[87][66], dotarray[88][66], dotarray[89][66], dotarray[90][66], dotarray[91][66], dotarray[92][66], dotarray[93][66], dotarray[94][66], dotarray[95][66], dotarray[96][66], dotarray[97][66], dotarray[98][66], dotarray[99][66], dotarray[100][66], dotarray[101][66], dotarray[102][66], dotarray[103][66], dotarray[104][66], dotarray[105][66], dotarray[106][66], dotarray[107][66], dotarray[108][66], dotarray[109][66], dotarray[110][66], dotarray[111][66], dotarray[112][66], dotarray[113][66], dotarray[114][66], dotarray[115][66], dotarray[116][66], dotarray[117][66], dotarray[118][66], dotarray[119][66], dotarray[120][66], dotarray[121][66], dotarray[122][66], dotarray[123][66], dotarray[124][66], dotarray[125][66], dotarray[126][66], dotarray[127][66]};
assign dot_col_67 = {dotarray[0][67], dotarray[1][67], dotarray[2][67], dotarray[3][67], dotarray[4][67], dotarray[5][67], dotarray[6][67], dotarray[7][67], dotarray[8][67], dotarray[9][67], dotarray[10][67], dotarray[11][67], dotarray[12][67], dotarray[13][67], dotarray[14][67], dotarray[15][67], dotarray[16][67], dotarray[17][67], dotarray[18][67], dotarray[19][67], dotarray[20][67], dotarray[21][67], dotarray[22][67], dotarray[23][67], dotarray[24][67], dotarray[25][67], dotarray[26][67], dotarray[27][67], dotarray[28][67], dotarray[29][67], dotarray[30][67], dotarray[31][67], dotarray[32][67], dotarray[33][67], dotarray[34][67], dotarray[35][67], dotarray[36][67], dotarray[37][67], dotarray[38][67], dotarray[39][67], dotarray[40][67], dotarray[41][67], dotarray[42][67], dotarray[43][67], dotarray[44][67], dotarray[45][67], dotarray[46][67], dotarray[47][67], dotarray[48][67], dotarray[49][67], dotarray[50][67], dotarray[51][67], dotarray[52][67], dotarray[53][67], dotarray[54][67], dotarray[55][67], dotarray[56][67], dotarray[57][67], dotarray[58][67], dotarray[59][67], dotarray[60][67], dotarray[61][67], dotarray[62][67], dotarray[63][67], dotarray[64][67], dotarray[65][67], dotarray[66][67], dotarray[67][67], dotarray[68][67], dotarray[69][67], dotarray[70][67], dotarray[71][67], dotarray[72][67], dotarray[73][67], dotarray[74][67], dotarray[75][67], dotarray[76][67], dotarray[77][67], dotarray[78][67], dotarray[79][67], dotarray[80][67], dotarray[81][67], dotarray[82][67], dotarray[83][67], dotarray[84][67], dotarray[85][67], dotarray[86][67], dotarray[87][67], dotarray[88][67], dotarray[89][67], dotarray[90][67], dotarray[91][67], dotarray[92][67], dotarray[93][67], dotarray[94][67], dotarray[95][67], dotarray[96][67], dotarray[97][67], dotarray[98][67], dotarray[99][67], dotarray[100][67], dotarray[101][67], dotarray[102][67], dotarray[103][67], dotarray[104][67], dotarray[105][67], dotarray[106][67], dotarray[107][67], dotarray[108][67], dotarray[109][67], dotarray[110][67], dotarray[111][67], dotarray[112][67], dotarray[113][67], dotarray[114][67], dotarray[115][67], dotarray[116][67], dotarray[117][67], dotarray[118][67], dotarray[119][67], dotarray[120][67], dotarray[121][67], dotarray[122][67], dotarray[123][67], dotarray[124][67], dotarray[125][67], dotarray[126][67], dotarray[127][67]};
assign dot_col_68 = {dotarray[0][68], dotarray[1][68], dotarray[2][68], dotarray[3][68], dotarray[4][68], dotarray[5][68], dotarray[6][68], dotarray[7][68], dotarray[8][68], dotarray[9][68], dotarray[10][68], dotarray[11][68], dotarray[12][68], dotarray[13][68], dotarray[14][68], dotarray[15][68], dotarray[16][68], dotarray[17][68], dotarray[18][68], dotarray[19][68], dotarray[20][68], dotarray[21][68], dotarray[22][68], dotarray[23][68], dotarray[24][68], dotarray[25][68], dotarray[26][68], dotarray[27][68], dotarray[28][68], dotarray[29][68], dotarray[30][68], dotarray[31][68], dotarray[32][68], dotarray[33][68], dotarray[34][68], dotarray[35][68], dotarray[36][68], dotarray[37][68], dotarray[38][68], dotarray[39][68], dotarray[40][68], dotarray[41][68], dotarray[42][68], dotarray[43][68], dotarray[44][68], dotarray[45][68], dotarray[46][68], dotarray[47][68], dotarray[48][68], dotarray[49][68], dotarray[50][68], dotarray[51][68], dotarray[52][68], dotarray[53][68], dotarray[54][68], dotarray[55][68], dotarray[56][68], dotarray[57][68], dotarray[58][68], dotarray[59][68], dotarray[60][68], dotarray[61][68], dotarray[62][68], dotarray[63][68], dotarray[64][68], dotarray[65][68], dotarray[66][68], dotarray[67][68], dotarray[68][68], dotarray[69][68], dotarray[70][68], dotarray[71][68], dotarray[72][68], dotarray[73][68], dotarray[74][68], dotarray[75][68], dotarray[76][68], dotarray[77][68], dotarray[78][68], dotarray[79][68], dotarray[80][68], dotarray[81][68], dotarray[82][68], dotarray[83][68], dotarray[84][68], dotarray[85][68], dotarray[86][68], dotarray[87][68], dotarray[88][68], dotarray[89][68], dotarray[90][68], dotarray[91][68], dotarray[92][68], dotarray[93][68], dotarray[94][68], dotarray[95][68], dotarray[96][68], dotarray[97][68], dotarray[98][68], dotarray[99][68], dotarray[100][68], dotarray[101][68], dotarray[102][68], dotarray[103][68], dotarray[104][68], dotarray[105][68], dotarray[106][68], dotarray[107][68], dotarray[108][68], dotarray[109][68], dotarray[110][68], dotarray[111][68], dotarray[112][68], dotarray[113][68], dotarray[114][68], dotarray[115][68], dotarray[116][68], dotarray[117][68], dotarray[118][68], dotarray[119][68], dotarray[120][68], dotarray[121][68], dotarray[122][68], dotarray[123][68], dotarray[124][68], dotarray[125][68], dotarray[126][68], dotarray[127][68]};
assign dot_col_69 = {dotarray[0][69], dotarray[1][69], dotarray[2][69], dotarray[3][69], dotarray[4][69], dotarray[5][69], dotarray[6][69], dotarray[7][69], dotarray[8][69], dotarray[9][69], dotarray[10][69], dotarray[11][69], dotarray[12][69], dotarray[13][69], dotarray[14][69], dotarray[15][69], dotarray[16][69], dotarray[17][69], dotarray[18][69], dotarray[19][69], dotarray[20][69], dotarray[21][69], dotarray[22][69], dotarray[23][69], dotarray[24][69], dotarray[25][69], dotarray[26][69], dotarray[27][69], dotarray[28][69], dotarray[29][69], dotarray[30][69], dotarray[31][69], dotarray[32][69], dotarray[33][69], dotarray[34][69], dotarray[35][69], dotarray[36][69], dotarray[37][69], dotarray[38][69], dotarray[39][69], dotarray[40][69], dotarray[41][69], dotarray[42][69], dotarray[43][69], dotarray[44][69], dotarray[45][69], dotarray[46][69], dotarray[47][69], dotarray[48][69], dotarray[49][69], dotarray[50][69], dotarray[51][69], dotarray[52][69], dotarray[53][69], dotarray[54][69], dotarray[55][69], dotarray[56][69], dotarray[57][69], dotarray[58][69], dotarray[59][69], dotarray[60][69], dotarray[61][69], dotarray[62][69], dotarray[63][69], dotarray[64][69], dotarray[65][69], dotarray[66][69], dotarray[67][69], dotarray[68][69], dotarray[69][69], dotarray[70][69], dotarray[71][69], dotarray[72][69], dotarray[73][69], dotarray[74][69], dotarray[75][69], dotarray[76][69], dotarray[77][69], dotarray[78][69], dotarray[79][69], dotarray[80][69], dotarray[81][69], dotarray[82][69], dotarray[83][69], dotarray[84][69], dotarray[85][69], dotarray[86][69], dotarray[87][69], dotarray[88][69], dotarray[89][69], dotarray[90][69], dotarray[91][69], dotarray[92][69], dotarray[93][69], dotarray[94][69], dotarray[95][69], dotarray[96][69], dotarray[97][69], dotarray[98][69], dotarray[99][69], dotarray[100][69], dotarray[101][69], dotarray[102][69], dotarray[103][69], dotarray[104][69], dotarray[105][69], dotarray[106][69], dotarray[107][69], dotarray[108][69], dotarray[109][69], dotarray[110][69], dotarray[111][69], dotarray[112][69], dotarray[113][69], dotarray[114][69], dotarray[115][69], dotarray[116][69], dotarray[117][69], dotarray[118][69], dotarray[119][69], dotarray[120][69], dotarray[121][69], dotarray[122][69], dotarray[123][69], dotarray[124][69], dotarray[125][69], dotarray[126][69], dotarray[127][69]};
assign dot_col_70 = {dotarray[0][70], dotarray[1][70], dotarray[2][70], dotarray[3][70], dotarray[4][70], dotarray[5][70], dotarray[6][70], dotarray[7][70], dotarray[8][70], dotarray[9][70], dotarray[10][70], dotarray[11][70], dotarray[12][70], dotarray[13][70], dotarray[14][70], dotarray[15][70], dotarray[16][70], dotarray[17][70], dotarray[18][70], dotarray[19][70], dotarray[20][70], dotarray[21][70], dotarray[22][70], dotarray[23][70], dotarray[24][70], dotarray[25][70], dotarray[26][70], dotarray[27][70], dotarray[28][70], dotarray[29][70], dotarray[30][70], dotarray[31][70], dotarray[32][70], dotarray[33][70], dotarray[34][70], dotarray[35][70], dotarray[36][70], dotarray[37][70], dotarray[38][70], dotarray[39][70], dotarray[40][70], dotarray[41][70], dotarray[42][70], dotarray[43][70], dotarray[44][70], dotarray[45][70], dotarray[46][70], dotarray[47][70], dotarray[48][70], dotarray[49][70], dotarray[50][70], dotarray[51][70], dotarray[52][70], dotarray[53][70], dotarray[54][70], dotarray[55][70], dotarray[56][70], dotarray[57][70], dotarray[58][70], dotarray[59][70], dotarray[60][70], dotarray[61][70], dotarray[62][70], dotarray[63][70], dotarray[64][70], dotarray[65][70], dotarray[66][70], dotarray[67][70], dotarray[68][70], dotarray[69][70], dotarray[70][70], dotarray[71][70], dotarray[72][70], dotarray[73][70], dotarray[74][70], dotarray[75][70], dotarray[76][70], dotarray[77][70], dotarray[78][70], dotarray[79][70], dotarray[80][70], dotarray[81][70], dotarray[82][70], dotarray[83][70], dotarray[84][70], dotarray[85][70], dotarray[86][70], dotarray[87][70], dotarray[88][70], dotarray[89][70], dotarray[90][70], dotarray[91][70], dotarray[92][70], dotarray[93][70], dotarray[94][70], dotarray[95][70], dotarray[96][70], dotarray[97][70], dotarray[98][70], dotarray[99][70], dotarray[100][70], dotarray[101][70], dotarray[102][70], dotarray[103][70], dotarray[104][70], dotarray[105][70], dotarray[106][70], dotarray[107][70], dotarray[108][70], dotarray[109][70], dotarray[110][70], dotarray[111][70], dotarray[112][70], dotarray[113][70], dotarray[114][70], dotarray[115][70], dotarray[116][70], dotarray[117][70], dotarray[118][70], dotarray[119][70], dotarray[120][70], dotarray[121][70], dotarray[122][70], dotarray[123][70], dotarray[124][70], dotarray[125][70], dotarray[126][70], dotarray[127][70]};
assign dot_col_71 = {dotarray[0][71], dotarray[1][71], dotarray[2][71], dotarray[3][71], dotarray[4][71], dotarray[5][71], dotarray[6][71], dotarray[7][71], dotarray[8][71], dotarray[9][71], dotarray[10][71], dotarray[11][71], dotarray[12][71], dotarray[13][71], dotarray[14][71], dotarray[15][71], dotarray[16][71], dotarray[17][71], dotarray[18][71], dotarray[19][71], dotarray[20][71], dotarray[21][71], dotarray[22][71], dotarray[23][71], dotarray[24][71], dotarray[25][71], dotarray[26][71], dotarray[27][71], dotarray[28][71], dotarray[29][71], dotarray[30][71], dotarray[31][71], dotarray[32][71], dotarray[33][71], dotarray[34][71], dotarray[35][71], dotarray[36][71], dotarray[37][71], dotarray[38][71], dotarray[39][71], dotarray[40][71], dotarray[41][71], dotarray[42][71], dotarray[43][71], dotarray[44][71], dotarray[45][71], dotarray[46][71], dotarray[47][71], dotarray[48][71], dotarray[49][71], dotarray[50][71], dotarray[51][71], dotarray[52][71], dotarray[53][71], dotarray[54][71], dotarray[55][71], dotarray[56][71], dotarray[57][71], dotarray[58][71], dotarray[59][71], dotarray[60][71], dotarray[61][71], dotarray[62][71], dotarray[63][71], dotarray[64][71], dotarray[65][71], dotarray[66][71], dotarray[67][71], dotarray[68][71], dotarray[69][71], dotarray[70][71], dotarray[71][71], dotarray[72][71], dotarray[73][71], dotarray[74][71], dotarray[75][71], dotarray[76][71], dotarray[77][71], dotarray[78][71], dotarray[79][71], dotarray[80][71], dotarray[81][71], dotarray[82][71], dotarray[83][71], dotarray[84][71], dotarray[85][71], dotarray[86][71], dotarray[87][71], dotarray[88][71], dotarray[89][71], dotarray[90][71], dotarray[91][71], dotarray[92][71], dotarray[93][71], dotarray[94][71], dotarray[95][71], dotarray[96][71], dotarray[97][71], dotarray[98][71], dotarray[99][71], dotarray[100][71], dotarray[101][71], dotarray[102][71], dotarray[103][71], dotarray[104][71], dotarray[105][71], dotarray[106][71], dotarray[107][71], dotarray[108][71], dotarray[109][71], dotarray[110][71], dotarray[111][71], dotarray[112][71], dotarray[113][71], dotarray[114][71], dotarray[115][71], dotarray[116][71], dotarray[117][71], dotarray[118][71], dotarray[119][71], dotarray[120][71], dotarray[121][71], dotarray[122][71], dotarray[123][71], dotarray[124][71], dotarray[125][71], dotarray[126][71], dotarray[127][71]};
assign dot_col_72 = {dotarray[0][72], dotarray[1][72], dotarray[2][72], dotarray[3][72], dotarray[4][72], dotarray[5][72], dotarray[6][72], dotarray[7][72], dotarray[8][72], dotarray[9][72], dotarray[10][72], dotarray[11][72], dotarray[12][72], dotarray[13][72], dotarray[14][72], dotarray[15][72], dotarray[16][72], dotarray[17][72], dotarray[18][72], dotarray[19][72], dotarray[20][72], dotarray[21][72], dotarray[22][72], dotarray[23][72], dotarray[24][72], dotarray[25][72], dotarray[26][72], dotarray[27][72], dotarray[28][72], dotarray[29][72], dotarray[30][72], dotarray[31][72], dotarray[32][72], dotarray[33][72], dotarray[34][72], dotarray[35][72], dotarray[36][72], dotarray[37][72], dotarray[38][72], dotarray[39][72], dotarray[40][72], dotarray[41][72], dotarray[42][72], dotarray[43][72], dotarray[44][72], dotarray[45][72], dotarray[46][72], dotarray[47][72], dotarray[48][72], dotarray[49][72], dotarray[50][72], dotarray[51][72], dotarray[52][72], dotarray[53][72], dotarray[54][72], dotarray[55][72], dotarray[56][72], dotarray[57][72], dotarray[58][72], dotarray[59][72], dotarray[60][72], dotarray[61][72], dotarray[62][72], dotarray[63][72], dotarray[64][72], dotarray[65][72], dotarray[66][72], dotarray[67][72], dotarray[68][72], dotarray[69][72], dotarray[70][72], dotarray[71][72], dotarray[72][72], dotarray[73][72], dotarray[74][72], dotarray[75][72], dotarray[76][72], dotarray[77][72], dotarray[78][72], dotarray[79][72], dotarray[80][72], dotarray[81][72], dotarray[82][72], dotarray[83][72], dotarray[84][72], dotarray[85][72], dotarray[86][72], dotarray[87][72], dotarray[88][72], dotarray[89][72], dotarray[90][72], dotarray[91][72], dotarray[92][72], dotarray[93][72], dotarray[94][72], dotarray[95][72], dotarray[96][72], dotarray[97][72], dotarray[98][72], dotarray[99][72], dotarray[100][72], dotarray[101][72], dotarray[102][72], dotarray[103][72], dotarray[104][72], dotarray[105][72], dotarray[106][72], dotarray[107][72], dotarray[108][72], dotarray[109][72], dotarray[110][72], dotarray[111][72], dotarray[112][72], dotarray[113][72], dotarray[114][72], dotarray[115][72], dotarray[116][72], dotarray[117][72], dotarray[118][72], dotarray[119][72], dotarray[120][72], dotarray[121][72], dotarray[122][72], dotarray[123][72], dotarray[124][72], dotarray[125][72], dotarray[126][72], dotarray[127][72]};
assign dot_col_73 = {dotarray[0][73], dotarray[1][73], dotarray[2][73], dotarray[3][73], dotarray[4][73], dotarray[5][73], dotarray[6][73], dotarray[7][73], dotarray[8][73], dotarray[9][73], dotarray[10][73], dotarray[11][73], dotarray[12][73], dotarray[13][73], dotarray[14][73], dotarray[15][73], dotarray[16][73], dotarray[17][73], dotarray[18][73], dotarray[19][73], dotarray[20][73], dotarray[21][73], dotarray[22][73], dotarray[23][73], dotarray[24][73], dotarray[25][73], dotarray[26][73], dotarray[27][73], dotarray[28][73], dotarray[29][73], dotarray[30][73], dotarray[31][73], dotarray[32][73], dotarray[33][73], dotarray[34][73], dotarray[35][73], dotarray[36][73], dotarray[37][73], dotarray[38][73], dotarray[39][73], dotarray[40][73], dotarray[41][73], dotarray[42][73], dotarray[43][73], dotarray[44][73], dotarray[45][73], dotarray[46][73], dotarray[47][73], dotarray[48][73], dotarray[49][73], dotarray[50][73], dotarray[51][73], dotarray[52][73], dotarray[53][73], dotarray[54][73], dotarray[55][73], dotarray[56][73], dotarray[57][73], dotarray[58][73], dotarray[59][73], dotarray[60][73], dotarray[61][73], dotarray[62][73], dotarray[63][73], dotarray[64][73], dotarray[65][73], dotarray[66][73], dotarray[67][73], dotarray[68][73], dotarray[69][73], dotarray[70][73], dotarray[71][73], dotarray[72][73], dotarray[73][73], dotarray[74][73], dotarray[75][73], dotarray[76][73], dotarray[77][73], dotarray[78][73], dotarray[79][73], dotarray[80][73], dotarray[81][73], dotarray[82][73], dotarray[83][73], dotarray[84][73], dotarray[85][73], dotarray[86][73], dotarray[87][73], dotarray[88][73], dotarray[89][73], dotarray[90][73], dotarray[91][73], dotarray[92][73], dotarray[93][73], dotarray[94][73], dotarray[95][73], dotarray[96][73], dotarray[97][73], dotarray[98][73], dotarray[99][73], dotarray[100][73], dotarray[101][73], dotarray[102][73], dotarray[103][73], dotarray[104][73], dotarray[105][73], dotarray[106][73], dotarray[107][73], dotarray[108][73], dotarray[109][73], dotarray[110][73], dotarray[111][73], dotarray[112][73], dotarray[113][73], dotarray[114][73], dotarray[115][73], dotarray[116][73], dotarray[117][73], dotarray[118][73], dotarray[119][73], dotarray[120][73], dotarray[121][73], dotarray[122][73], dotarray[123][73], dotarray[124][73], dotarray[125][73], dotarray[126][73], dotarray[127][73]};
assign dot_col_74 = {dotarray[0][74], dotarray[1][74], dotarray[2][74], dotarray[3][74], dotarray[4][74], dotarray[5][74], dotarray[6][74], dotarray[7][74], dotarray[8][74], dotarray[9][74], dotarray[10][74], dotarray[11][74], dotarray[12][74], dotarray[13][74], dotarray[14][74], dotarray[15][74], dotarray[16][74], dotarray[17][74], dotarray[18][74], dotarray[19][74], dotarray[20][74], dotarray[21][74], dotarray[22][74], dotarray[23][74], dotarray[24][74], dotarray[25][74], dotarray[26][74], dotarray[27][74], dotarray[28][74], dotarray[29][74], dotarray[30][74], dotarray[31][74], dotarray[32][74], dotarray[33][74], dotarray[34][74], dotarray[35][74], dotarray[36][74], dotarray[37][74], dotarray[38][74], dotarray[39][74], dotarray[40][74], dotarray[41][74], dotarray[42][74], dotarray[43][74], dotarray[44][74], dotarray[45][74], dotarray[46][74], dotarray[47][74], dotarray[48][74], dotarray[49][74], dotarray[50][74], dotarray[51][74], dotarray[52][74], dotarray[53][74], dotarray[54][74], dotarray[55][74], dotarray[56][74], dotarray[57][74], dotarray[58][74], dotarray[59][74], dotarray[60][74], dotarray[61][74], dotarray[62][74], dotarray[63][74], dotarray[64][74], dotarray[65][74], dotarray[66][74], dotarray[67][74], dotarray[68][74], dotarray[69][74], dotarray[70][74], dotarray[71][74], dotarray[72][74], dotarray[73][74], dotarray[74][74], dotarray[75][74], dotarray[76][74], dotarray[77][74], dotarray[78][74], dotarray[79][74], dotarray[80][74], dotarray[81][74], dotarray[82][74], dotarray[83][74], dotarray[84][74], dotarray[85][74], dotarray[86][74], dotarray[87][74], dotarray[88][74], dotarray[89][74], dotarray[90][74], dotarray[91][74], dotarray[92][74], dotarray[93][74], dotarray[94][74], dotarray[95][74], dotarray[96][74], dotarray[97][74], dotarray[98][74], dotarray[99][74], dotarray[100][74], dotarray[101][74], dotarray[102][74], dotarray[103][74], dotarray[104][74], dotarray[105][74], dotarray[106][74], dotarray[107][74], dotarray[108][74], dotarray[109][74], dotarray[110][74], dotarray[111][74], dotarray[112][74], dotarray[113][74], dotarray[114][74], dotarray[115][74], dotarray[116][74], dotarray[117][74], dotarray[118][74], dotarray[119][74], dotarray[120][74], dotarray[121][74], dotarray[122][74], dotarray[123][74], dotarray[124][74], dotarray[125][74], dotarray[126][74], dotarray[127][74]};
assign dot_col_75 = {dotarray[0][75], dotarray[1][75], dotarray[2][75], dotarray[3][75], dotarray[4][75], dotarray[5][75], dotarray[6][75], dotarray[7][75], dotarray[8][75], dotarray[9][75], dotarray[10][75], dotarray[11][75], dotarray[12][75], dotarray[13][75], dotarray[14][75], dotarray[15][75], dotarray[16][75], dotarray[17][75], dotarray[18][75], dotarray[19][75], dotarray[20][75], dotarray[21][75], dotarray[22][75], dotarray[23][75], dotarray[24][75], dotarray[25][75], dotarray[26][75], dotarray[27][75], dotarray[28][75], dotarray[29][75], dotarray[30][75], dotarray[31][75], dotarray[32][75], dotarray[33][75], dotarray[34][75], dotarray[35][75], dotarray[36][75], dotarray[37][75], dotarray[38][75], dotarray[39][75], dotarray[40][75], dotarray[41][75], dotarray[42][75], dotarray[43][75], dotarray[44][75], dotarray[45][75], dotarray[46][75], dotarray[47][75], dotarray[48][75], dotarray[49][75], dotarray[50][75], dotarray[51][75], dotarray[52][75], dotarray[53][75], dotarray[54][75], dotarray[55][75], dotarray[56][75], dotarray[57][75], dotarray[58][75], dotarray[59][75], dotarray[60][75], dotarray[61][75], dotarray[62][75], dotarray[63][75], dotarray[64][75], dotarray[65][75], dotarray[66][75], dotarray[67][75], dotarray[68][75], dotarray[69][75], dotarray[70][75], dotarray[71][75], dotarray[72][75], dotarray[73][75], dotarray[74][75], dotarray[75][75], dotarray[76][75], dotarray[77][75], dotarray[78][75], dotarray[79][75], dotarray[80][75], dotarray[81][75], dotarray[82][75], dotarray[83][75], dotarray[84][75], dotarray[85][75], dotarray[86][75], dotarray[87][75], dotarray[88][75], dotarray[89][75], dotarray[90][75], dotarray[91][75], dotarray[92][75], dotarray[93][75], dotarray[94][75], dotarray[95][75], dotarray[96][75], dotarray[97][75], dotarray[98][75], dotarray[99][75], dotarray[100][75], dotarray[101][75], dotarray[102][75], dotarray[103][75], dotarray[104][75], dotarray[105][75], dotarray[106][75], dotarray[107][75], dotarray[108][75], dotarray[109][75], dotarray[110][75], dotarray[111][75], dotarray[112][75], dotarray[113][75], dotarray[114][75], dotarray[115][75], dotarray[116][75], dotarray[117][75], dotarray[118][75], dotarray[119][75], dotarray[120][75], dotarray[121][75], dotarray[122][75], dotarray[123][75], dotarray[124][75], dotarray[125][75], dotarray[126][75], dotarray[127][75]};
assign dot_col_76 = {dotarray[0][76], dotarray[1][76], dotarray[2][76], dotarray[3][76], dotarray[4][76], dotarray[5][76], dotarray[6][76], dotarray[7][76], dotarray[8][76], dotarray[9][76], dotarray[10][76], dotarray[11][76], dotarray[12][76], dotarray[13][76], dotarray[14][76], dotarray[15][76], dotarray[16][76], dotarray[17][76], dotarray[18][76], dotarray[19][76], dotarray[20][76], dotarray[21][76], dotarray[22][76], dotarray[23][76], dotarray[24][76], dotarray[25][76], dotarray[26][76], dotarray[27][76], dotarray[28][76], dotarray[29][76], dotarray[30][76], dotarray[31][76], dotarray[32][76], dotarray[33][76], dotarray[34][76], dotarray[35][76], dotarray[36][76], dotarray[37][76], dotarray[38][76], dotarray[39][76], dotarray[40][76], dotarray[41][76], dotarray[42][76], dotarray[43][76], dotarray[44][76], dotarray[45][76], dotarray[46][76], dotarray[47][76], dotarray[48][76], dotarray[49][76], dotarray[50][76], dotarray[51][76], dotarray[52][76], dotarray[53][76], dotarray[54][76], dotarray[55][76], dotarray[56][76], dotarray[57][76], dotarray[58][76], dotarray[59][76], dotarray[60][76], dotarray[61][76], dotarray[62][76], dotarray[63][76], dotarray[64][76], dotarray[65][76], dotarray[66][76], dotarray[67][76], dotarray[68][76], dotarray[69][76], dotarray[70][76], dotarray[71][76], dotarray[72][76], dotarray[73][76], dotarray[74][76], dotarray[75][76], dotarray[76][76], dotarray[77][76], dotarray[78][76], dotarray[79][76], dotarray[80][76], dotarray[81][76], dotarray[82][76], dotarray[83][76], dotarray[84][76], dotarray[85][76], dotarray[86][76], dotarray[87][76], dotarray[88][76], dotarray[89][76], dotarray[90][76], dotarray[91][76], dotarray[92][76], dotarray[93][76], dotarray[94][76], dotarray[95][76], dotarray[96][76], dotarray[97][76], dotarray[98][76], dotarray[99][76], dotarray[100][76], dotarray[101][76], dotarray[102][76], dotarray[103][76], dotarray[104][76], dotarray[105][76], dotarray[106][76], dotarray[107][76], dotarray[108][76], dotarray[109][76], dotarray[110][76], dotarray[111][76], dotarray[112][76], dotarray[113][76], dotarray[114][76], dotarray[115][76], dotarray[116][76], dotarray[117][76], dotarray[118][76], dotarray[119][76], dotarray[120][76], dotarray[121][76], dotarray[122][76], dotarray[123][76], dotarray[124][76], dotarray[125][76], dotarray[126][76], dotarray[127][76]};
assign dot_col_77 = {dotarray[0][77], dotarray[1][77], dotarray[2][77], dotarray[3][77], dotarray[4][77], dotarray[5][77], dotarray[6][77], dotarray[7][77], dotarray[8][77], dotarray[9][77], dotarray[10][77], dotarray[11][77], dotarray[12][77], dotarray[13][77], dotarray[14][77], dotarray[15][77], dotarray[16][77], dotarray[17][77], dotarray[18][77], dotarray[19][77], dotarray[20][77], dotarray[21][77], dotarray[22][77], dotarray[23][77], dotarray[24][77], dotarray[25][77], dotarray[26][77], dotarray[27][77], dotarray[28][77], dotarray[29][77], dotarray[30][77], dotarray[31][77], dotarray[32][77], dotarray[33][77], dotarray[34][77], dotarray[35][77], dotarray[36][77], dotarray[37][77], dotarray[38][77], dotarray[39][77], dotarray[40][77], dotarray[41][77], dotarray[42][77], dotarray[43][77], dotarray[44][77], dotarray[45][77], dotarray[46][77], dotarray[47][77], dotarray[48][77], dotarray[49][77], dotarray[50][77], dotarray[51][77], dotarray[52][77], dotarray[53][77], dotarray[54][77], dotarray[55][77], dotarray[56][77], dotarray[57][77], dotarray[58][77], dotarray[59][77], dotarray[60][77], dotarray[61][77], dotarray[62][77], dotarray[63][77], dotarray[64][77], dotarray[65][77], dotarray[66][77], dotarray[67][77], dotarray[68][77], dotarray[69][77], dotarray[70][77], dotarray[71][77], dotarray[72][77], dotarray[73][77], dotarray[74][77], dotarray[75][77], dotarray[76][77], dotarray[77][77], dotarray[78][77], dotarray[79][77], dotarray[80][77], dotarray[81][77], dotarray[82][77], dotarray[83][77], dotarray[84][77], dotarray[85][77], dotarray[86][77], dotarray[87][77], dotarray[88][77], dotarray[89][77], dotarray[90][77], dotarray[91][77], dotarray[92][77], dotarray[93][77], dotarray[94][77], dotarray[95][77], dotarray[96][77], dotarray[97][77], dotarray[98][77], dotarray[99][77], dotarray[100][77], dotarray[101][77], dotarray[102][77], dotarray[103][77], dotarray[104][77], dotarray[105][77], dotarray[106][77], dotarray[107][77], dotarray[108][77], dotarray[109][77], dotarray[110][77], dotarray[111][77], dotarray[112][77], dotarray[113][77], dotarray[114][77], dotarray[115][77], dotarray[116][77], dotarray[117][77], dotarray[118][77], dotarray[119][77], dotarray[120][77], dotarray[121][77], dotarray[122][77], dotarray[123][77], dotarray[124][77], dotarray[125][77], dotarray[126][77], dotarray[127][77]};
assign dot_col_78 = {dotarray[0][78], dotarray[1][78], dotarray[2][78], dotarray[3][78], dotarray[4][78], dotarray[5][78], dotarray[6][78], dotarray[7][78], dotarray[8][78], dotarray[9][78], dotarray[10][78], dotarray[11][78], dotarray[12][78], dotarray[13][78], dotarray[14][78], dotarray[15][78], dotarray[16][78], dotarray[17][78], dotarray[18][78], dotarray[19][78], dotarray[20][78], dotarray[21][78], dotarray[22][78], dotarray[23][78], dotarray[24][78], dotarray[25][78], dotarray[26][78], dotarray[27][78], dotarray[28][78], dotarray[29][78], dotarray[30][78], dotarray[31][78], dotarray[32][78], dotarray[33][78], dotarray[34][78], dotarray[35][78], dotarray[36][78], dotarray[37][78], dotarray[38][78], dotarray[39][78], dotarray[40][78], dotarray[41][78], dotarray[42][78], dotarray[43][78], dotarray[44][78], dotarray[45][78], dotarray[46][78], dotarray[47][78], dotarray[48][78], dotarray[49][78], dotarray[50][78], dotarray[51][78], dotarray[52][78], dotarray[53][78], dotarray[54][78], dotarray[55][78], dotarray[56][78], dotarray[57][78], dotarray[58][78], dotarray[59][78], dotarray[60][78], dotarray[61][78], dotarray[62][78], dotarray[63][78], dotarray[64][78], dotarray[65][78], dotarray[66][78], dotarray[67][78], dotarray[68][78], dotarray[69][78], dotarray[70][78], dotarray[71][78], dotarray[72][78], dotarray[73][78], dotarray[74][78], dotarray[75][78], dotarray[76][78], dotarray[77][78], dotarray[78][78], dotarray[79][78], dotarray[80][78], dotarray[81][78], dotarray[82][78], dotarray[83][78], dotarray[84][78], dotarray[85][78], dotarray[86][78], dotarray[87][78], dotarray[88][78], dotarray[89][78], dotarray[90][78], dotarray[91][78], dotarray[92][78], dotarray[93][78], dotarray[94][78], dotarray[95][78], dotarray[96][78], dotarray[97][78], dotarray[98][78], dotarray[99][78], dotarray[100][78], dotarray[101][78], dotarray[102][78], dotarray[103][78], dotarray[104][78], dotarray[105][78], dotarray[106][78], dotarray[107][78], dotarray[108][78], dotarray[109][78], dotarray[110][78], dotarray[111][78], dotarray[112][78], dotarray[113][78], dotarray[114][78], dotarray[115][78], dotarray[116][78], dotarray[117][78], dotarray[118][78], dotarray[119][78], dotarray[120][78], dotarray[121][78], dotarray[122][78], dotarray[123][78], dotarray[124][78], dotarray[125][78], dotarray[126][78], dotarray[127][78]};
assign dot_col_79 = {dotarray[0][79], dotarray[1][79], dotarray[2][79], dotarray[3][79], dotarray[4][79], dotarray[5][79], dotarray[6][79], dotarray[7][79], dotarray[8][79], dotarray[9][79], dotarray[10][79], dotarray[11][79], dotarray[12][79], dotarray[13][79], dotarray[14][79], dotarray[15][79], dotarray[16][79], dotarray[17][79], dotarray[18][79], dotarray[19][79], dotarray[20][79], dotarray[21][79], dotarray[22][79], dotarray[23][79], dotarray[24][79], dotarray[25][79], dotarray[26][79], dotarray[27][79], dotarray[28][79], dotarray[29][79], dotarray[30][79], dotarray[31][79], dotarray[32][79], dotarray[33][79], dotarray[34][79], dotarray[35][79], dotarray[36][79], dotarray[37][79], dotarray[38][79], dotarray[39][79], dotarray[40][79], dotarray[41][79], dotarray[42][79], dotarray[43][79], dotarray[44][79], dotarray[45][79], dotarray[46][79], dotarray[47][79], dotarray[48][79], dotarray[49][79], dotarray[50][79], dotarray[51][79], dotarray[52][79], dotarray[53][79], dotarray[54][79], dotarray[55][79], dotarray[56][79], dotarray[57][79], dotarray[58][79], dotarray[59][79], dotarray[60][79], dotarray[61][79], dotarray[62][79], dotarray[63][79], dotarray[64][79], dotarray[65][79], dotarray[66][79], dotarray[67][79], dotarray[68][79], dotarray[69][79], dotarray[70][79], dotarray[71][79], dotarray[72][79], dotarray[73][79], dotarray[74][79], dotarray[75][79], dotarray[76][79], dotarray[77][79], dotarray[78][79], dotarray[79][79], dotarray[80][79], dotarray[81][79], dotarray[82][79], dotarray[83][79], dotarray[84][79], dotarray[85][79], dotarray[86][79], dotarray[87][79], dotarray[88][79], dotarray[89][79], dotarray[90][79], dotarray[91][79], dotarray[92][79], dotarray[93][79], dotarray[94][79], dotarray[95][79], dotarray[96][79], dotarray[97][79], dotarray[98][79], dotarray[99][79], dotarray[100][79], dotarray[101][79], dotarray[102][79], dotarray[103][79], dotarray[104][79], dotarray[105][79], dotarray[106][79], dotarray[107][79], dotarray[108][79], dotarray[109][79], dotarray[110][79], dotarray[111][79], dotarray[112][79], dotarray[113][79], dotarray[114][79], dotarray[115][79], dotarray[116][79], dotarray[117][79], dotarray[118][79], dotarray[119][79], dotarray[120][79], dotarray[121][79], dotarray[122][79], dotarray[123][79], dotarray[124][79], dotarray[125][79], dotarray[126][79], dotarray[127][79]};
assign dot_col_80 = {dotarray[0][80], dotarray[1][80], dotarray[2][80], dotarray[3][80], dotarray[4][80], dotarray[5][80], dotarray[6][80], dotarray[7][80], dotarray[8][80], dotarray[9][80], dotarray[10][80], dotarray[11][80], dotarray[12][80], dotarray[13][80], dotarray[14][80], dotarray[15][80], dotarray[16][80], dotarray[17][80], dotarray[18][80], dotarray[19][80], dotarray[20][80], dotarray[21][80], dotarray[22][80], dotarray[23][80], dotarray[24][80], dotarray[25][80], dotarray[26][80], dotarray[27][80], dotarray[28][80], dotarray[29][80], dotarray[30][80], dotarray[31][80], dotarray[32][80], dotarray[33][80], dotarray[34][80], dotarray[35][80], dotarray[36][80], dotarray[37][80], dotarray[38][80], dotarray[39][80], dotarray[40][80], dotarray[41][80], dotarray[42][80], dotarray[43][80], dotarray[44][80], dotarray[45][80], dotarray[46][80], dotarray[47][80], dotarray[48][80], dotarray[49][80], dotarray[50][80], dotarray[51][80], dotarray[52][80], dotarray[53][80], dotarray[54][80], dotarray[55][80], dotarray[56][80], dotarray[57][80], dotarray[58][80], dotarray[59][80], dotarray[60][80], dotarray[61][80], dotarray[62][80], dotarray[63][80], dotarray[64][80], dotarray[65][80], dotarray[66][80], dotarray[67][80], dotarray[68][80], dotarray[69][80], dotarray[70][80], dotarray[71][80], dotarray[72][80], dotarray[73][80], dotarray[74][80], dotarray[75][80], dotarray[76][80], dotarray[77][80], dotarray[78][80], dotarray[79][80], dotarray[80][80], dotarray[81][80], dotarray[82][80], dotarray[83][80], dotarray[84][80], dotarray[85][80], dotarray[86][80], dotarray[87][80], dotarray[88][80], dotarray[89][80], dotarray[90][80], dotarray[91][80], dotarray[92][80], dotarray[93][80], dotarray[94][80], dotarray[95][80], dotarray[96][80], dotarray[97][80], dotarray[98][80], dotarray[99][80], dotarray[100][80], dotarray[101][80], dotarray[102][80], dotarray[103][80], dotarray[104][80], dotarray[105][80], dotarray[106][80], dotarray[107][80], dotarray[108][80], dotarray[109][80], dotarray[110][80], dotarray[111][80], dotarray[112][80], dotarray[113][80], dotarray[114][80], dotarray[115][80], dotarray[116][80], dotarray[117][80], dotarray[118][80], dotarray[119][80], dotarray[120][80], dotarray[121][80], dotarray[122][80], dotarray[123][80], dotarray[124][80], dotarray[125][80], dotarray[126][80], dotarray[127][80]};
assign dot_col_81 = {dotarray[0][81], dotarray[1][81], dotarray[2][81], dotarray[3][81], dotarray[4][81], dotarray[5][81], dotarray[6][81], dotarray[7][81], dotarray[8][81], dotarray[9][81], dotarray[10][81], dotarray[11][81], dotarray[12][81], dotarray[13][81], dotarray[14][81], dotarray[15][81], dotarray[16][81], dotarray[17][81], dotarray[18][81], dotarray[19][81], dotarray[20][81], dotarray[21][81], dotarray[22][81], dotarray[23][81], dotarray[24][81], dotarray[25][81], dotarray[26][81], dotarray[27][81], dotarray[28][81], dotarray[29][81], dotarray[30][81], dotarray[31][81], dotarray[32][81], dotarray[33][81], dotarray[34][81], dotarray[35][81], dotarray[36][81], dotarray[37][81], dotarray[38][81], dotarray[39][81], dotarray[40][81], dotarray[41][81], dotarray[42][81], dotarray[43][81], dotarray[44][81], dotarray[45][81], dotarray[46][81], dotarray[47][81], dotarray[48][81], dotarray[49][81], dotarray[50][81], dotarray[51][81], dotarray[52][81], dotarray[53][81], dotarray[54][81], dotarray[55][81], dotarray[56][81], dotarray[57][81], dotarray[58][81], dotarray[59][81], dotarray[60][81], dotarray[61][81], dotarray[62][81], dotarray[63][81], dotarray[64][81], dotarray[65][81], dotarray[66][81], dotarray[67][81], dotarray[68][81], dotarray[69][81], dotarray[70][81], dotarray[71][81], dotarray[72][81], dotarray[73][81], dotarray[74][81], dotarray[75][81], dotarray[76][81], dotarray[77][81], dotarray[78][81], dotarray[79][81], dotarray[80][81], dotarray[81][81], dotarray[82][81], dotarray[83][81], dotarray[84][81], dotarray[85][81], dotarray[86][81], dotarray[87][81], dotarray[88][81], dotarray[89][81], dotarray[90][81], dotarray[91][81], dotarray[92][81], dotarray[93][81], dotarray[94][81], dotarray[95][81], dotarray[96][81], dotarray[97][81], dotarray[98][81], dotarray[99][81], dotarray[100][81], dotarray[101][81], dotarray[102][81], dotarray[103][81], dotarray[104][81], dotarray[105][81], dotarray[106][81], dotarray[107][81], dotarray[108][81], dotarray[109][81], dotarray[110][81], dotarray[111][81], dotarray[112][81], dotarray[113][81], dotarray[114][81], dotarray[115][81], dotarray[116][81], dotarray[117][81], dotarray[118][81], dotarray[119][81], dotarray[120][81], dotarray[121][81], dotarray[122][81], dotarray[123][81], dotarray[124][81], dotarray[125][81], dotarray[126][81], dotarray[127][81]};
assign dot_col_82 = {dotarray[0][82], dotarray[1][82], dotarray[2][82], dotarray[3][82], dotarray[4][82], dotarray[5][82], dotarray[6][82], dotarray[7][82], dotarray[8][82], dotarray[9][82], dotarray[10][82], dotarray[11][82], dotarray[12][82], dotarray[13][82], dotarray[14][82], dotarray[15][82], dotarray[16][82], dotarray[17][82], dotarray[18][82], dotarray[19][82], dotarray[20][82], dotarray[21][82], dotarray[22][82], dotarray[23][82], dotarray[24][82], dotarray[25][82], dotarray[26][82], dotarray[27][82], dotarray[28][82], dotarray[29][82], dotarray[30][82], dotarray[31][82], dotarray[32][82], dotarray[33][82], dotarray[34][82], dotarray[35][82], dotarray[36][82], dotarray[37][82], dotarray[38][82], dotarray[39][82], dotarray[40][82], dotarray[41][82], dotarray[42][82], dotarray[43][82], dotarray[44][82], dotarray[45][82], dotarray[46][82], dotarray[47][82], dotarray[48][82], dotarray[49][82], dotarray[50][82], dotarray[51][82], dotarray[52][82], dotarray[53][82], dotarray[54][82], dotarray[55][82], dotarray[56][82], dotarray[57][82], dotarray[58][82], dotarray[59][82], dotarray[60][82], dotarray[61][82], dotarray[62][82], dotarray[63][82], dotarray[64][82], dotarray[65][82], dotarray[66][82], dotarray[67][82], dotarray[68][82], dotarray[69][82], dotarray[70][82], dotarray[71][82], dotarray[72][82], dotarray[73][82], dotarray[74][82], dotarray[75][82], dotarray[76][82], dotarray[77][82], dotarray[78][82], dotarray[79][82], dotarray[80][82], dotarray[81][82], dotarray[82][82], dotarray[83][82], dotarray[84][82], dotarray[85][82], dotarray[86][82], dotarray[87][82], dotarray[88][82], dotarray[89][82], dotarray[90][82], dotarray[91][82], dotarray[92][82], dotarray[93][82], dotarray[94][82], dotarray[95][82], dotarray[96][82], dotarray[97][82], dotarray[98][82], dotarray[99][82], dotarray[100][82], dotarray[101][82], dotarray[102][82], dotarray[103][82], dotarray[104][82], dotarray[105][82], dotarray[106][82], dotarray[107][82], dotarray[108][82], dotarray[109][82], dotarray[110][82], dotarray[111][82], dotarray[112][82], dotarray[113][82], dotarray[114][82], dotarray[115][82], dotarray[116][82], dotarray[117][82], dotarray[118][82], dotarray[119][82], dotarray[120][82], dotarray[121][82], dotarray[122][82], dotarray[123][82], dotarray[124][82], dotarray[125][82], dotarray[126][82], dotarray[127][82]};
assign dot_col_83 = {dotarray[0][83], dotarray[1][83], dotarray[2][83], dotarray[3][83], dotarray[4][83], dotarray[5][83], dotarray[6][83], dotarray[7][83], dotarray[8][83], dotarray[9][83], dotarray[10][83], dotarray[11][83], dotarray[12][83], dotarray[13][83], dotarray[14][83], dotarray[15][83], dotarray[16][83], dotarray[17][83], dotarray[18][83], dotarray[19][83], dotarray[20][83], dotarray[21][83], dotarray[22][83], dotarray[23][83], dotarray[24][83], dotarray[25][83], dotarray[26][83], dotarray[27][83], dotarray[28][83], dotarray[29][83], dotarray[30][83], dotarray[31][83], dotarray[32][83], dotarray[33][83], dotarray[34][83], dotarray[35][83], dotarray[36][83], dotarray[37][83], dotarray[38][83], dotarray[39][83], dotarray[40][83], dotarray[41][83], dotarray[42][83], dotarray[43][83], dotarray[44][83], dotarray[45][83], dotarray[46][83], dotarray[47][83], dotarray[48][83], dotarray[49][83], dotarray[50][83], dotarray[51][83], dotarray[52][83], dotarray[53][83], dotarray[54][83], dotarray[55][83], dotarray[56][83], dotarray[57][83], dotarray[58][83], dotarray[59][83], dotarray[60][83], dotarray[61][83], dotarray[62][83], dotarray[63][83], dotarray[64][83], dotarray[65][83], dotarray[66][83], dotarray[67][83], dotarray[68][83], dotarray[69][83], dotarray[70][83], dotarray[71][83], dotarray[72][83], dotarray[73][83], dotarray[74][83], dotarray[75][83], dotarray[76][83], dotarray[77][83], dotarray[78][83], dotarray[79][83], dotarray[80][83], dotarray[81][83], dotarray[82][83], dotarray[83][83], dotarray[84][83], dotarray[85][83], dotarray[86][83], dotarray[87][83], dotarray[88][83], dotarray[89][83], dotarray[90][83], dotarray[91][83], dotarray[92][83], dotarray[93][83], dotarray[94][83], dotarray[95][83], dotarray[96][83], dotarray[97][83], dotarray[98][83], dotarray[99][83], dotarray[100][83], dotarray[101][83], dotarray[102][83], dotarray[103][83], dotarray[104][83], dotarray[105][83], dotarray[106][83], dotarray[107][83], dotarray[108][83], dotarray[109][83], dotarray[110][83], dotarray[111][83], dotarray[112][83], dotarray[113][83], dotarray[114][83], dotarray[115][83], dotarray[116][83], dotarray[117][83], dotarray[118][83], dotarray[119][83], dotarray[120][83], dotarray[121][83], dotarray[122][83], dotarray[123][83], dotarray[124][83], dotarray[125][83], dotarray[126][83], dotarray[127][83]};
assign dot_col_84 = {dotarray[0][84], dotarray[1][84], dotarray[2][84], dotarray[3][84], dotarray[4][84], dotarray[5][84], dotarray[6][84], dotarray[7][84], dotarray[8][84], dotarray[9][84], dotarray[10][84], dotarray[11][84], dotarray[12][84], dotarray[13][84], dotarray[14][84], dotarray[15][84], dotarray[16][84], dotarray[17][84], dotarray[18][84], dotarray[19][84], dotarray[20][84], dotarray[21][84], dotarray[22][84], dotarray[23][84], dotarray[24][84], dotarray[25][84], dotarray[26][84], dotarray[27][84], dotarray[28][84], dotarray[29][84], dotarray[30][84], dotarray[31][84], dotarray[32][84], dotarray[33][84], dotarray[34][84], dotarray[35][84], dotarray[36][84], dotarray[37][84], dotarray[38][84], dotarray[39][84], dotarray[40][84], dotarray[41][84], dotarray[42][84], dotarray[43][84], dotarray[44][84], dotarray[45][84], dotarray[46][84], dotarray[47][84], dotarray[48][84], dotarray[49][84], dotarray[50][84], dotarray[51][84], dotarray[52][84], dotarray[53][84], dotarray[54][84], dotarray[55][84], dotarray[56][84], dotarray[57][84], dotarray[58][84], dotarray[59][84], dotarray[60][84], dotarray[61][84], dotarray[62][84], dotarray[63][84], dotarray[64][84], dotarray[65][84], dotarray[66][84], dotarray[67][84], dotarray[68][84], dotarray[69][84], dotarray[70][84], dotarray[71][84], dotarray[72][84], dotarray[73][84], dotarray[74][84], dotarray[75][84], dotarray[76][84], dotarray[77][84], dotarray[78][84], dotarray[79][84], dotarray[80][84], dotarray[81][84], dotarray[82][84], dotarray[83][84], dotarray[84][84], dotarray[85][84], dotarray[86][84], dotarray[87][84], dotarray[88][84], dotarray[89][84], dotarray[90][84], dotarray[91][84], dotarray[92][84], dotarray[93][84], dotarray[94][84], dotarray[95][84], dotarray[96][84], dotarray[97][84], dotarray[98][84], dotarray[99][84], dotarray[100][84], dotarray[101][84], dotarray[102][84], dotarray[103][84], dotarray[104][84], dotarray[105][84], dotarray[106][84], dotarray[107][84], dotarray[108][84], dotarray[109][84], dotarray[110][84], dotarray[111][84], dotarray[112][84], dotarray[113][84], dotarray[114][84], dotarray[115][84], dotarray[116][84], dotarray[117][84], dotarray[118][84], dotarray[119][84], dotarray[120][84], dotarray[121][84], dotarray[122][84], dotarray[123][84], dotarray[124][84], dotarray[125][84], dotarray[126][84], dotarray[127][84]};
assign dot_col_85 = {dotarray[0][85], dotarray[1][85], dotarray[2][85], dotarray[3][85], dotarray[4][85], dotarray[5][85], dotarray[6][85], dotarray[7][85], dotarray[8][85], dotarray[9][85], dotarray[10][85], dotarray[11][85], dotarray[12][85], dotarray[13][85], dotarray[14][85], dotarray[15][85], dotarray[16][85], dotarray[17][85], dotarray[18][85], dotarray[19][85], dotarray[20][85], dotarray[21][85], dotarray[22][85], dotarray[23][85], dotarray[24][85], dotarray[25][85], dotarray[26][85], dotarray[27][85], dotarray[28][85], dotarray[29][85], dotarray[30][85], dotarray[31][85], dotarray[32][85], dotarray[33][85], dotarray[34][85], dotarray[35][85], dotarray[36][85], dotarray[37][85], dotarray[38][85], dotarray[39][85], dotarray[40][85], dotarray[41][85], dotarray[42][85], dotarray[43][85], dotarray[44][85], dotarray[45][85], dotarray[46][85], dotarray[47][85], dotarray[48][85], dotarray[49][85], dotarray[50][85], dotarray[51][85], dotarray[52][85], dotarray[53][85], dotarray[54][85], dotarray[55][85], dotarray[56][85], dotarray[57][85], dotarray[58][85], dotarray[59][85], dotarray[60][85], dotarray[61][85], dotarray[62][85], dotarray[63][85], dotarray[64][85], dotarray[65][85], dotarray[66][85], dotarray[67][85], dotarray[68][85], dotarray[69][85], dotarray[70][85], dotarray[71][85], dotarray[72][85], dotarray[73][85], dotarray[74][85], dotarray[75][85], dotarray[76][85], dotarray[77][85], dotarray[78][85], dotarray[79][85], dotarray[80][85], dotarray[81][85], dotarray[82][85], dotarray[83][85], dotarray[84][85], dotarray[85][85], dotarray[86][85], dotarray[87][85], dotarray[88][85], dotarray[89][85], dotarray[90][85], dotarray[91][85], dotarray[92][85], dotarray[93][85], dotarray[94][85], dotarray[95][85], dotarray[96][85], dotarray[97][85], dotarray[98][85], dotarray[99][85], dotarray[100][85], dotarray[101][85], dotarray[102][85], dotarray[103][85], dotarray[104][85], dotarray[105][85], dotarray[106][85], dotarray[107][85], dotarray[108][85], dotarray[109][85], dotarray[110][85], dotarray[111][85], dotarray[112][85], dotarray[113][85], dotarray[114][85], dotarray[115][85], dotarray[116][85], dotarray[117][85], dotarray[118][85], dotarray[119][85], dotarray[120][85], dotarray[121][85], dotarray[122][85], dotarray[123][85], dotarray[124][85], dotarray[125][85], dotarray[126][85], dotarray[127][85]};
assign dot_col_86 = {dotarray[0][86], dotarray[1][86], dotarray[2][86], dotarray[3][86], dotarray[4][86], dotarray[5][86], dotarray[6][86], dotarray[7][86], dotarray[8][86], dotarray[9][86], dotarray[10][86], dotarray[11][86], dotarray[12][86], dotarray[13][86], dotarray[14][86], dotarray[15][86], dotarray[16][86], dotarray[17][86], dotarray[18][86], dotarray[19][86], dotarray[20][86], dotarray[21][86], dotarray[22][86], dotarray[23][86], dotarray[24][86], dotarray[25][86], dotarray[26][86], dotarray[27][86], dotarray[28][86], dotarray[29][86], dotarray[30][86], dotarray[31][86], dotarray[32][86], dotarray[33][86], dotarray[34][86], dotarray[35][86], dotarray[36][86], dotarray[37][86], dotarray[38][86], dotarray[39][86], dotarray[40][86], dotarray[41][86], dotarray[42][86], dotarray[43][86], dotarray[44][86], dotarray[45][86], dotarray[46][86], dotarray[47][86], dotarray[48][86], dotarray[49][86], dotarray[50][86], dotarray[51][86], dotarray[52][86], dotarray[53][86], dotarray[54][86], dotarray[55][86], dotarray[56][86], dotarray[57][86], dotarray[58][86], dotarray[59][86], dotarray[60][86], dotarray[61][86], dotarray[62][86], dotarray[63][86], dotarray[64][86], dotarray[65][86], dotarray[66][86], dotarray[67][86], dotarray[68][86], dotarray[69][86], dotarray[70][86], dotarray[71][86], dotarray[72][86], dotarray[73][86], dotarray[74][86], dotarray[75][86], dotarray[76][86], dotarray[77][86], dotarray[78][86], dotarray[79][86], dotarray[80][86], dotarray[81][86], dotarray[82][86], dotarray[83][86], dotarray[84][86], dotarray[85][86], dotarray[86][86], dotarray[87][86], dotarray[88][86], dotarray[89][86], dotarray[90][86], dotarray[91][86], dotarray[92][86], dotarray[93][86], dotarray[94][86], dotarray[95][86], dotarray[96][86], dotarray[97][86], dotarray[98][86], dotarray[99][86], dotarray[100][86], dotarray[101][86], dotarray[102][86], dotarray[103][86], dotarray[104][86], dotarray[105][86], dotarray[106][86], dotarray[107][86], dotarray[108][86], dotarray[109][86], dotarray[110][86], dotarray[111][86], dotarray[112][86], dotarray[113][86], dotarray[114][86], dotarray[115][86], dotarray[116][86], dotarray[117][86], dotarray[118][86], dotarray[119][86], dotarray[120][86], dotarray[121][86], dotarray[122][86], dotarray[123][86], dotarray[124][86], dotarray[125][86], dotarray[126][86], dotarray[127][86]};
assign dot_col_87 = {dotarray[0][87], dotarray[1][87], dotarray[2][87], dotarray[3][87], dotarray[4][87], dotarray[5][87], dotarray[6][87], dotarray[7][87], dotarray[8][87], dotarray[9][87], dotarray[10][87], dotarray[11][87], dotarray[12][87], dotarray[13][87], dotarray[14][87], dotarray[15][87], dotarray[16][87], dotarray[17][87], dotarray[18][87], dotarray[19][87], dotarray[20][87], dotarray[21][87], dotarray[22][87], dotarray[23][87], dotarray[24][87], dotarray[25][87], dotarray[26][87], dotarray[27][87], dotarray[28][87], dotarray[29][87], dotarray[30][87], dotarray[31][87], dotarray[32][87], dotarray[33][87], dotarray[34][87], dotarray[35][87], dotarray[36][87], dotarray[37][87], dotarray[38][87], dotarray[39][87], dotarray[40][87], dotarray[41][87], dotarray[42][87], dotarray[43][87], dotarray[44][87], dotarray[45][87], dotarray[46][87], dotarray[47][87], dotarray[48][87], dotarray[49][87], dotarray[50][87], dotarray[51][87], dotarray[52][87], dotarray[53][87], dotarray[54][87], dotarray[55][87], dotarray[56][87], dotarray[57][87], dotarray[58][87], dotarray[59][87], dotarray[60][87], dotarray[61][87], dotarray[62][87], dotarray[63][87], dotarray[64][87], dotarray[65][87], dotarray[66][87], dotarray[67][87], dotarray[68][87], dotarray[69][87], dotarray[70][87], dotarray[71][87], dotarray[72][87], dotarray[73][87], dotarray[74][87], dotarray[75][87], dotarray[76][87], dotarray[77][87], dotarray[78][87], dotarray[79][87], dotarray[80][87], dotarray[81][87], dotarray[82][87], dotarray[83][87], dotarray[84][87], dotarray[85][87], dotarray[86][87], dotarray[87][87], dotarray[88][87], dotarray[89][87], dotarray[90][87], dotarray[91][87], dotarray[92][87], dotarray[93][87], dotarray[94][87], dotarray[95][87], dotarray[96][87], dotarray[97][87], dotarray[98][87], dotarray[99][87], dotarray[100][87], dotarray[101][87], dotarray[102][87], dotarray[103][87], dotarray[104][87], dotarray[105][87], dotarray[106][87], dotarray[107][87], dotarray[108][87], dotarray[109][87], dotarray[110][87], dotarray[111][87], dotarray[112][87], dotarray[113][87], dotarray[114][87], dotarray[115][87], dotarray[116][87], dotarray[117][87], dotarray[118][87], dotarray[119][87], dotarray[120][87], dotarray[121][87], dotarray[122][87], dotarray[123][87], dotarray[124][87], dotarray[125][87], dotarray[126][87], dotarray[127][87]};
assign dot_col_88 = {dotarray[0][88], dotarray[1][88], dotarray[2][88], dotarray[3][88], dotarray[4][88], dotarray[5][88], dotarray[6][88], dotarray[7][88], dotarray[8][88], dotarray[9][88], dotarray[10][88], dotarray[11][88], dotarray[12][88], dotarray[13][88], dotarray[14][88], dotarray[15][88], dotarray[16][88], dotarray[17][88], dotarray[18][88], dotarray[19][88], dotarray[20][88], dotarray[21][88], dotarray[22][88], dotarray[23][88], dotarray[24][88], dotarray[25][88], dotarray[26][88], dotarray[27][88], dotarray[28][88], dotarray[29][88], dotarray[30][88], dotarray[31][88], dotarray[32][88], dotarray[33][88], dotarray[34][88], dotarray[35][88], dotarray[36][88], dotarray[37][88], dotarray[38][88], dotarray[39][88], dotarray[40][88], dotarray[41][88], dotarray[42][88], dotarray[43][88], dotarray[44][88], dotarray[45][88], dotarray[46][88], dotarray[47][88], dotarray[48][88], dotarray[49][88], dotarray[50][88], dotarray[51][88], dotarray[52][88], dotarray[53][88], dotarray[54][88], dotarray[55][88], dotarray[56][88], dotarray[57][88], dotarray[58][88], dotarray[59][88], dotarray[60][88], dotarray[61][88], dotarray[62][88], dotarray[63][88], dotarray[64][88], dotarray[65][88], dotarray[66][88], dotarray[67][88], dotarray[68][88], dotarray[69][88], dotarray[70][88], dotarray[71][88], dotarray[72][88], dotarray[73][88], dotarray[74][88], dotarray[75][88], dotarray[76][88], dotarray[77][88], dotarray[78][88], dotarray[79][88], dotarray[80][88], dotarray[81][88], dotarray[82][88], dotarray[83][88], dotarray[84][88], dotarray[85][88], dotarray[86][88], dotarray[87][88], dotarray[88][88], dotarray[89][88], dotarray[90][88], dotarray[91][88], dotarray[92][88], dotarray[93][88], dotarray[94][88], dotarray[95][88], dotarray[96][88], dotarray[97][88], dotarray[98][88], dotarray[99][88], dotarray[100][88], dotarray[101][88], dotarray[102][88], dotarray[103][88], dotarray[104][88], dotarray[105][88], dotarray[106][88], dotarray[107][88], dotarray[108][88], dotarray[109][88], dotarray[110][88], dotarray[111][88], dotarray[112][88], dotarray[113][88], dotarray[114][88], dotarray[115][88], dotarray[116][88], dotarray[117][88], dotarray[118][88], dotarray[119][88], dotarray[120][88], dotarray[121][88], dotarray[122][88], dotarray[123][88], dotarray[124][88], dotarray[125][88], dotarray[126][88], dotarray[127][88]};
assign dot_col_89 = {dotarray[0][89], dotarray[1][89], dotarray[2][89], dotarray[3][89], dotarray[4][89], dotarray[5][89], dotarray[6][89], dotarray[7][89], dotarray[8][89], dotarray[9][89], dotarray[10][89], dotarray[11][89], dotarray[12][89], dotarray[13][89], dotarray[14][89], dotarray[15][89], dotarray[16][89], dotarray[17][89], dotarray[18][89], dotarray[19][89], dotarray[20][89], dotarray[21][89], dotarray[22][89], dotarray[23][89], dotarray[24][89], dotarray[25][89], dotarray[26][89], dotarray[27][89], dotarray[28][89], dotarray[29][89], dotarray[30][89], dotarray[31][89], dotarray[32][89], dotarray[33][89], dotarray[34][89], dotarray[35][89], dotarray[36][89], dotarray[37][89], dotarray[38][89], dotarray[39][89], dotarray[40][89], dotarray[41][89], dotarray[42][89], dotarray[43][89], dotarray[44][89], dotarray[45][89], dotarray[46][89], dotarray[47][89], dotarray[48][89], dotarray[49][89], dotarray[50][89], dotarray[51][89], dotarray[52][89], dotarray[53][89], dotarray[54][89], dotarray[55][89], dotarray[56][89], dotarray[57][89], dotarray[58][89], dotarray[59][89], dotarray[60][89], dotarray[61][89], dotarray[62][89], dotarray[63][89], dotarray[64][89], dotarray[65][89], dotarray[66][89], dotarray[67][89], dotarray[68][89], dotarray[69][89], dotarray[70][89], dotarray[71][89], dotarray[72][89], dotarray[73][89], dotarray[74][89], dotarray[75][89], dotarray[76][89], dotarray[77][89], dotarray[78][89], dotarray[79][89], dotarray[80][89], dotarray[81][89], dotarray[82][89], dotarray[83][89], dotarray[84][89], dotarray[85][89], dotarray[86][89], dotarray[87][89], dotarray[88][89], dotarray[89][89], dotarray[90][89], dotarray[91][89], dotarray[92][89], dotarray[93][89], dotarray[94][89], dotarray[95][89], dotarray[96][89], dotarray[97][89], dotarray[98][89], dotarray[99][89], dotarray[100][89], dotarray[101][89], dotarray[102][89], dotarray[103][89], dotarray[104][89], dotarray[105][89], dotarray[106][89], dotarray[107][89], dotarray[108][89], dotarray[109][89], dotarray[110][89], dotarray[111][89], dotarray[112][89], dotarray[113][89], dotarray[114][89], dotarray[115][89], dotarray[116][89], dotarray[117][89], dotarray[118][89], dotarray[119][89], dotarray[120][89], dotarray[121][89], dotarray[122][89], dotarray[123][89], dotarray[124][89], dotarray[125][89], dotarray[126][89], dotarray[127][89]};
assign dot_col_90 = {dotarray[0][90], dotarray[1][90], dotarray[2][90], dotarray[3][90], dotarray[4][90], dotarray[5][90], dotarray[6][90], dotarray[7][90], dotarray[8][90], dotarray[9][90], dotarray[10][90], dotarray[11][90], dotarray[12][90], dotarray[13][90], dotarray[14][90], dotarray[15][90], dotarray[16][90], dotarray[17][90], dotarray[18][90], dotarray[19][90], dotarray[20][90], dotarray[21][90], dotarray[22][90], dotarray[23][90], dotarray[24][90], dotarray[25][90], dotarray[26][90], dotarray[27][90], dotarray[28][90], dotarray[29][90], dotarray[30][90], dotarray[31][90], dotarray[32][90], dotarray[33][90], dotarray[34][90], dotarray[35][90], dotarray[36][90], dotarray[37][90], dotarray[38][90], dotarray[39][90], dotarray[40][90], dotarray[41][90], dotarray[42][90], dotarray[43][90], dotarray[44][90], dotarray[45][90], dotarray[46][90], dotarray[47][90], dotarray[48][90], dotarray[49][90], dotarray[50][90], dotarray[51][90], dotarray[52][90], dotarray[53][90], dotarray[54][90], dotarray[55][90], dotarray[56][90], dotarray[57][90], dotarray[58][90], dotarray[59][90], dotarray[60][90], dotarray[61][90], dotarray[62][90], dotarray[63][90], dotarray[64][90], dotarray[65][90], dotarray[66][90], dotarray[67][90], dotarray[68][90], dotarray[69][90], dotarray[70][90], dotarray[71][90], dotarray[72][90], dotarray[73][90], dotarray[74][90], dotarray[75][90], dotarray[76][90], dotarray[77][90], dotarray[78][90], dotarray[79][90], dotarray[80][90], dotarray[81][90], dotarray[82][90], dotarray[83][90], dotarray[84][90], dotarray[85][90], dotarray[86][90], dotarray[87][90], dotarray[88][90], dotarray[89][90], dotarray[90][90], dotarray[91][90], dotarray[92][90], dotarray[93][90], dotarray[94][90], dotarray[95][90], dotarray[96][90], dotarray[97][90], dotarray[98][90], dotarray[99][90], dotarray[100][90], dotarray[101][90], dotarray[102][90], dotarray[103][90], dotarray[104][90], dotarray[105][90], dotarray[106][90], dotarray[107][90], dotarray[108][90], dotarray[109][90], dotarray[110][90], dotarray[111][90], dotarray[112][90], dotarray[113][90], dotarray[114][90], dotarray[115][90], dotarray[116][90], dotarray[117][90], dotarray[118][90], dotarray[119][90], dotarray[120][90], dotarray[121][90], dotarray[122][90], dotarray[123][90], dotarray[124][90], dotarray[125][90], dotarray[126][90], dotarray[127][90]};
assign dot_col_91 = {dotarray[0][91], dotarray[1][91], dotarray[2][91], dotarray[3][91], dotarray[4][91], dotarray[5][91], dotarray[6][91], dotarray[7][91], dotarray[8][91], dotarray[9][91], dotarray[10][91], dotarray[11][91], dotarray[12][91], dotarray[13][91], dotarray[14][91], dotarray[15][91], dotarray[16][91], dotarray[17][91], dotarray[18][91], dotarray[19][91], dotarray[20][91], dotarray[21][91], dotarray[22][91], dotarray[23][91], dotarray[24][91], dotarray[25][91], dotarray[26][91], dotarray[27][91], dotarray[28][91], dotarray[29][91], dotarray[30][91], dotarray[31][91], dotarray[32][91], dotarray[33][91], dotarray[34][91], dotarray[35][91], dotarray[36][91], dotarray[37][91], dotarray[38][91], dotarray[39][91], dotarray[40][91], dotarray[41][91], dotarray[42][91], dotarray[43][91], dotarray[44][91], dotarray[45][91], dotarray[46][91], dotarray[47][91], dotarray[48][91], dotarray[49][91], dotarray[50][91], dotarray[51][91], dotarray[52][91], dotarray[53][91], dotarray[54][91], dotarray[55][91], dotarray[56][91], dotarray[57][91], dotarray[58][91], dotarray[59][91], dotarray[60][91], dotarray[61][91], dotarray[62][91], dotarray[63][91], dotarray[64][91], dotarray[65][91], dotarray[66][91], dotarray[67][91], dotarray[68][91], dotarray[69][91], dotarray[70][91], dotarray[71][91], dotarray[72][91], dotarray[73][91], dotarray[74][91], dotarray[75][91], dotarray[76][91], dotarray[77][91], dotarray[78][91], dotarray[79][91], dotarray[80][91], dotarray[81][91], dotarray[82][91], dotarray[83][91], dotarray[84][91], dotarray[85][91], dotarray[86][91], dotarray[87][91], dotarray[88][91], dotarray[89][91], dotarray[90][91], dotarray[91][91], dotarray[92][91], dotarray[93][91], dotarray[94][91], dotarray[95][91], dotarray[96][91], dotarray[97][91], dotarray[98][91], dotarray[99][91], dotarray[100][91], dotarray[101][91], dotarray[102][91], dotarray[103][91], dotarray[104][91], dotarray[105][91], dotarray[106][91], dotarray[107][91], dotarray[108][91], dotarray[109][91], dotarray[110][91], dotarray[111][91], dotarray[112][91], dotarray[113][91], dotarray[114][91], dotarray[115][91], dotarray[116][91], dotarray[117][91], dotarray[118][91], dotarray[119][91], dotarray[120][91], dotarray[121][91], dotarray[122][91], dotarray[123][91], dotarray[124][91], dotarray[125][91], dotarray[126][91], dotarray[127][91]};
assign dot_col_92 = {dotarray[0][92], dotarray[1][92], dotarray[2][92], dotarray[3][92], dotarray[4][92], dotarray[5][92], dotarray[6][92], dotarray[7][92], dotarray[8][92], dotarray[9][92], dotarray[10][92], dotarray[11][92], dotarray[12][92], dotarray[13][92], dotarray[14][92], dotarray[15][92], dotarray[16][92], dotarray[17][92], dotarray[18][92], dotarray[19][92], dotarray[20][92], dotarray[21][92], dotarray[22][92], dotarray[23][92], dotarray[24][92], dotarray[25][92], dotarray[26][92], dotarray[27][92], dotarray[28][92], dotarray[29][92], dotarray[30][92], dotarray[31][92], dotarray[32][92], dotarray[33][92], dotarray[34][92], dotarray[35][92], dotarray[36][92], dotarray[37][92], dotarray[38][92], dotarray[39][92], dotarray[40][92], dotarray[41][92], dotarray[42][92], dotarray[43][92], dotarray[44][92], dotarray[45][92], dotarray[46][92], dotarray[47][92], dotarray[48][92], dotarray[49][92], dotarray[50][92], dotarray[51][92], dotarray[52][92], dotarray[53][92], dotarray[54][92], dotarray[55][92], dotarray[56][92], dotarray[57][92], dotarray[58][92], dotarray[59][92], dotarray[60][92], dotarray[61][92], dotarray[62][92], dotarray[63][92], dotarray[64][92], dotarray[65][92], dotarray[66][92], dotarray[67][92], dotarray[68][92], dotarray[69][92], dotarray[70][92], dotarray[71][92], dotarray[72][92], dotarray[73][92], dotarray[74][92], dotarray[75][92], dotarray[76][92], dotarray[77][92], dotarray[78][92], dotarray[79][92], dotarray[80][92], dotarray[81][92], dotarray[82][92], dotarray[83][92], dotarray[84][92], dotarray[85][92], dotarray[86][92], dotarray[87][92], dotarray[88][92], dotarray[89][92], dotarray[90][92], dotarray[91][92], dotarray[92][92], dotarray[93][92], dotarray[94][92], dotarray[95][92], dotarray[96][92], dotarray[97][92], dotarray[98][92], dotarray[99][92], dotarray[100][92], dotarray[101][92], dotarray[102][92], dotarray[103][92], dotarray[104][92], dotarray[105][92], dotarray[106][92], dotarray[107][92], dotarray[108][92], dotarray[109][92], dotarray[110][92], dotarray[111][92], dotarray[112][92], dotarray[113][92], dotarray[114][92], dotarray[115][92], dotarray[116][92], dotarray[117][92], dotarray[118][92], dotarray[119][92], dotarray[120][92], dotarray[121][92], dotarray[122][92], dotarray[123][92], dotarray[124][92], dotarray[125][92], dotarray[126][92], dotarray[127][92]};
assign dot_col_93 = {dotarray[0][93], dotarray[1][93], dotarray[2][93], dotarray[3][93], dotarray[4][93], dotarray[5][93], dotarray[6][93], dotarray[7][93], dotarray[8][93], dotarray[9][93], dotarray[10][93], dotarray[11][93], dotarray[12][93], dotarray[13][93], dotarray[14][93], dotarray[15][93], dotarray[16][93], dotarray[17][93], dotarray[18][93], dotarray[19][93], dotarray[20][93], dotarray[21][93], dotarray[22][93], dotarray[23][93], dotarray[24][93], dotarray[25][93], dotarray[26][93], dotarray[27][93], dotarray[28][93], dotarray[29][93], dotarray[30][93], dotarray[31][93], dotarray[32][93], dotarray[33][93], dotarray[34][93], dotarray[35][93], dotarray[36][93], dotarray[37][93], dotarray[38][93], dotarray[39][93], dotarray[40][93], dotarray[41][93], dotarray[42][93], dotarray[43][93], dotarray[44][93], dotarray[45][93], dotarray[46][93], dotarray[47][93], dotarray[48][93], dotarray[49][93], dotarray[50][93], dotarray[51][93], dotarray[52][93], dotarray[53][93], dotarray[54][93], dotarray[55][93], dotarray[56][93], dotarray[57][93], dotarray[58][93], dotarray[59][93], dotarray[60][93], dotarray[61][93], dotarray[62][93], dotarray[63][93], dotarray[64][93], dotarray[65][93], dotarray[66][93], dotarray[67][93], dotarray[68][93], dotarray[69][93], dotarray[70][93], dotarray[71][93], dotarray[72][93], dotarray[73][93], dotarray[74][93], dotarray[75][93], dotarray[76][93], dotarray[77][93], dotarray[78][93], dotarray[79][93], dotarray[80][93], dotarray[81][93], dotarray[82][93], dotarray[83][93], dotarray[84][93], dotarray[85][93], dotarray[86][93], dotarray[87][93], dotarray[88][93], dotarray[89][93], dotarray[90][93], dotarray[91][93], dotarray[92][93], dotarray[93][93], dotarray[94][93], dotarray[95][93], dotarray[96][93], dotarray[97][93], dotarray[98][93], dotarray[99][93], dotarray[100][93], dotarray[101][93], dotarray[102][93], dotarray[103][93], dotarray[104][93], dotarray[105][93], dotarray[106][93], dotarray[107][93], dotarray[108][93], dotarray[109][93], dotarray[110][93], dotarray[111][93], dotarray[112][93], dotarray[113][93], dotarray[114][93], dotarray[115][93], dotarray[116][93], dotarray[117][93], dotarray[118][93], dotarray[119][93], dotarray[120][93], dotarray[121][93], dotarray[122][93], dotarray[123][93], dotarray[124][93], dotarray[125][93], dotarray[126][93], dotarray[127][93]};
assign dot_col_94 = {dotarray[0][94], dotarray[1][94], dotarray[2][94], dotarray[3][94], dotarray[4][94], dotarray[5][94], dotarray[6][94], dotarray[7][94], dotarray[8][94], dotarray[9][94], dotarray[10][94], dotarray[11][94], dotarray[12][94], dotarray[13][94], dotarray[14][94], dotarray[15][94], dotarray[16][94], dotarray[17][94], dotarray[18][94], dotarray[19][94], dotarray[20][94], dotarray[21][94], dotarray[22][94], dotarray[23][94], dotarray[24][94], dotarray[25][94], dotarray[26][94], dotarray[27][94], dotarray[28][94], dotarray[29][94], dotarray[30][94], dotarray[31][94], dotarray[32][94], dotarray[33][94], dotarray[34][94], dotarray[35][94], dotarray[36][94], dotarray[37][94], dotarray[38][94], dotarray[39][94], dotarray[40][94], dotarray[41][94], dotarray[42][94], dotarray[43][94], dotarray[44][94], dotarray[45][94], dotarray[46][94], dotarray[47][94], dotarray[48][94], dotarray[49][94], dotarray[50][94], dotarray[51][94], dotarray[52][94], dotarray[53][94], dotarray[54][94], dotarray[55][94], dotarray[56][94], dotarray[57][94], dotarray[58][94], dotarray[59][94], dotarray[60][94], dotarray[61][94], dotarray[62][94], dotarray[63][94], dotarray[64][94], dotarray[65][94], dotarray[66][94], dotarray[67][94], dotarray[68][94], dotarray[69][94], dotarray[70][94], dotarray[71][94], dotarray[72][94], dotarray[73][94], dotarray[74][94], dotarray[75][94], dotarray[76][94], dotarray[77][94], dotarray[78][94], dotarray[79][94], dotarray[80][94], dotarray[81][94], dotarray[82][94], dotarray[83][94], dotarray[84][94], dotarray[85][94], dotarray[86][94], dotarray[87][94], dotarray[88][94], dotarray[89][94], dotarray[90][94], dotarray[91][94], dotarray[92][94], dotarray[93][94], dotarray[94][94], dotarray[95][94], dotarray[96][94], dotarray[97][94], dotarray[98][94], dotarray[99][94], dotarray[100][94], dotarray[101][94], dotarray[102][94], dotarray[103][94], dotarray[104][94], dotarray[105][94], dotarray[106][94], dotarray[107][94], dotarray[108][94], dotarray[109][94], dotarray[110][94], dotarray[111][94], dotarray[112][94], dotarray[113][94], dotarray[114][94], dotarray[115][94], dotarray[116][94], dotarray[117][94], dotarray[118][94], dotarray[119][94], dotarray[120][94], dotarray[121][94], dotarray[122][94], dotarray[123][94], dotarray[124][94], dotarray[125][94], dotarray[126][94], dotarray[127][94]};
assign dot_col_95 = {dotarray[0][95], dotarray[1][95], dotarray[2][95], dotarray[3][95], dotarray[4][95], dotarray[5][95], dotarray[6][95], dotarray[7][95], dotarray[8][95], dotarray[9][95], dotarray[10][95], dotarray[11][95], dotarray[12][95], dotarray[13][95], dotarray[14][95], dotarray[15][95], dotarray[16][95], dotarray[17][95], dotarray[18][95], dotarray[19][95], dotarray[20][95], dotarray[21][95], dotarray[22][95], dotarray[23][95], dotarray[24][95], dotarray[25][95], dotarray[26][95], dotarray[27][95], dotarray[28][95], dotarray[29][95], dotarray[30][95], dotarray[31][95], dotarray[32][95], dotarray[33][95], dotarray[34][95], dotarray[35][95], dotarray[36][95], dotarray[37][95], dotarray[38][95], dotarray[39][95], dotarray[40][95], dotarray[41][95], dotarray[42][95], dotarray[43][95], dotarray[44][95], dotarray[45][95], dotarray[46][95], dotarray[47][95], dotarray[48][95], dotarray[49][95], dotarray[50][95], dotarray[51][95], dotarray[52][95], dotarray[53][95], dotarray[54][95], dotarray[55][95], dotarray[56][95], dotarray[57][95], dotarray[58][95], dotarray[59][95], dotarray[60][95], dotarray[61][95], dotarray[62][95], dotarray[63][95], dotarray[64][95], dotarray[65][95], dotarray[66][95], dotarray[67][95], dotarray[68][95], dotarray[69][95], dotarray[70][95], dotarray[71][95], dotarray[72][95], dotarray[73][95], dotarray[74][95], dotarray[75][95], dotarray[76][95], dotarray[77][95], dotarray[78][95], dotarray[79][95], dotarray[80][95], dotarray[81][95], dotarray[82][95], dotarray[83][95], dotarray[84][95], dotarray[85][95], dotarray[86][95], dotarray[87][95], dotarray[88][95], dotarray[89][95], dotarray[90][95], dotarray[91][95], dotarray[92][95], dotarray[93][95], dotarray[94][95], dotarray[95][95], dotarray[96][95], dotarray[97][95], dotarray[98][95], dotarray[99][95], dotarray[100][95], dotarray[101][95], dotarray[102][95], dotarray[103][95], dotarray[104][95], dotarray[105][95], dotarray[106][95], dotarray[107][95], dotarray[108][95], dotarray[109][95], dotarray[110][95], dotarray[111][95], dotarray[112][95], dotarray[113][95], dotarray[114][95], dotarray[115][95], dotarray[116][95], dotarray[117][95], dotarray[118][95], dotarray[119][95], dotarray[120][95], dotarray[121][95], dotarray[122][95], dotarray[123][95], dotarray[124][95], dotarray[125][95], dotarray[126][95], dotarray[127][95]};
assign dot_col_96 = {dotarray[0][96], dotarray[1][96], dotarray[2][96], dotarray[3][96], dotarray[4][96], dotarray[5][96], dotarray[6][96], dotarray[7][96], dotarray[8][96], dotarray[9][96], dotarray[10][96], dotarray[11][96], dotarray[12][96], dotarray[13][96], dotarray[14][96], dotarray[15][96], dotarray[16][96], dotarray[17][96], dotarray[18][96], dotarray[19][96], dotarray[20][96], dotarray[21][96], dotarray[22][96], dotarray[23][96], dotarray[24][96], dotarray[25][96], dotarray[26][96], dotarray[27][96], dotarray[28][96], dotarray[29][96], dotarray[30][96], dotarray[31][96], dotarray[32][96], dotarray[33][96], dotarray[34][96], dotarray[35][96], dotarray[36][96], dotarray[37][96], dotarray[38][96], dotarray[39][96], dotarray[40][96], dotarray[41][96], dotarray[42][96], dotarray[43][96], dotarray[44][96], dotarray[45][96], dotarray[46][96], dotarray[47][96], dotarray[48][96], dotarray[49][96], dotarray[50][96], dotarray[51][96], dotarray[52][96], dotarray[53][96], dotarray[54][96], dotarray[55][96], dotarray[56][96], dotarray[57][96], dotarray[58][96], dotarray[59][96], dotarray[60][96], dotarray[61][96], dotarray[62][96], dotarray[63][96], dotarray[64][96], dotarray[65][96], dotarray[66][96], dotarray[67][96], dotarray[68][96], dotarray[69][96], dotarray[70][96], dotarray[71][96], dotarray[72][96], dotarray[73][96], dotarray[74][96], dotarray[75][96], dotarray[76][96], dotarray[77][96], dotarray[78][96], dotarray[79][96], dotarray[80][96], dotarray[81][96], dotarray[82][96], dotarray[83][96], dotarray[84][96], dotarray[85][96], dotarray[86][96], dotarray[87][96], dotarray[88][96], dotarray[89][96], dotarray[90][96], dotarray[91][96], dotarray[92][96], dotarray[93][96], dotarray[94][96], dotarray[95][96], dotarray[96][96], dotarray[97][96], dotarray[98][96], dotarray[99][96], dotarray[100][96], dotarray[101][96], dotarray[102][96], dotarray[103][96], dotarray[104][96], dotarray[105][96], dotarray[106][96], dotarray[107][96], dotarray[108][96], dotarray[109][96], dotarray[110][96], dotarray[111][96], dotarray[112][96], dotarray[113][96], dotarray[114][96], dotarray[115][96], dotarray[116][96], dotarray[117][96], dotarray[118][96], dotarray[119][96], dotarray[120][96], dotarray[121][96], dotarray[122][96], dotarray[123][96], dotarray[124][96], dotarray[125][96], dotarray[126][96], dotarray[127][96]};
assign dot_col_97 = {dotarray[0][97], dotarray[1][97], dotarray[2][97], dotarray[3][97], dotarray[4][97], dotarray[5][97], dotarray[6][97], dotarray[7][97], dotarray[8][97], dotarray[9][97], dotarray[10][97], dotarray[11][97], dotarray[12][97], dotarray[13][97], dotarray[14][97], dotarray[15][97], dotarray[16][97], dotarray[17][97], dotarray[18][97], dotarray[19][97], dotarray[20][97], dotarray[21][97], dotarray[22][97], dotarray[23][97], dotarray[24][97], dotarray[25][97], dotarray[26][97], dotarray[27][97], dotarray[28][97], dotarray[29][97], dotarray[30][97], dotarray[31][97], dotarray[32][97], dotarray[33][97], dotarray[34][97], dotarray[35][97], dotarray[36][97], dotarray[37][97], dotarray[38][97], dotarray[39][97], dotarray[40][97], dotarray[41][97], dotarray[42][97], dotarray[43][97], dotarray[44][97], dotarray[45][97], dotarray[46][97], dotarray[47][97], dotarray[48][97], dotarray[49][97], dotarray[50][97], dotarray[51][97], dotarray[52][97], dotarray[53][97], dotarray[54][97], dotarray[55][97], dotarray[56][97], dotarray[57][97], dotarray[58][97], dotarray[59][97], dotarray[60][97], dotarray[61][97], dotarray[62][97], dotarray[63][97], dotarray[64][97], dotarray[65][97], dotarray[66][97], dotarray[67][97], dotarray[68][97], dotarray[69][97], dotarray[70][97], dotarray[71][97], dotarray[72][97], dotarray[73][97], dotarray[74][97], dotarray[75][97], dotarray[76][97], dotarray[77][97], dotarray[78][97], dotarray[79][97], dotarray[80][97], dotarray[81][97], dotarray[82][97], dotarray[83][97], dotarray[84][97], dotarray[85][97], dotarray[86][97], dotarray[87][97], dotarray[88][97], dotarray[89][97], dotarray[90][97], dotarray[91][97], dotarray[92][97], dotarray[93][97], dotarray[94][97], dotarray[95][97], dotarray[96][97], dotarray[97][97], dotarray[98][97], dotarray[99][97], dotarray[100][97], dotarray[101][97], dotarray[102][97], dotarray[103][97], dotarray[104][97], dotarray[105][97], dotarray[106][97], dotarray[107][97], dotarray[108][97], dotarray[109][97], dotarray[110][97], dotarray[111][97], dotarray[112][97], dotarray[113][97], dotarray[114][97], dotarray[115][97], dotarray[116][97], dotarray[117][97], dotarray[118][97], dotarray[119][97], dotarray[120][97], dotarray[121][97], dotarray[122][97], dotarray[123][97], dotarray[124][97], dotarray[125][97], dotarray[126][97], dotarray[127][97]};
assign dot_col_98 = {dotarray[0][98], dotarray[1][98], dotarray[2][98], dotarray[3][98], dotarray[4][98], dotarray[5][98], dotarray[6][98], dotarray[7][98], dotarray[8][98], dotarray[9][98], dotarray[10][98], dotarray[11][98], dotarray[12][98], dotarray[13][98], dotarray[14][98], dotarray[15][98], dotarray[16][98], dotarray[17][98], dotarray[18][98], dotarray[19][98], dotarray[20][98], dotarray[21][98], dotarray[22][98], dotarray[23][98], dotarray[24][98], dotarray[25][98], dotarray[26][98], dotarray[27][98], dotarray[28][98], dotarray[29][98], dotarray[30][98], dotarray[31][98], dotarray[32][98], dotarray[33][98], dotarray[34][98], dotarray[35][98], dotarray[36][98], dotarray[37][98], dotarray[38][98], dotarray[39][98], dotarray[40][98], dotarray[41][98], dotarray[42][98], dotarray[43][98], dotarray[44][98], dotarray[45][98], dotarray[46][98], dotarray[47][98], dotarray[48][98], dotarray[49][98], dotarray[50][98], dotarray[51][98], dotarray[52][98], dotarray[53][98], dotarray[54][98], dotarray[55][98], dotarray[56][98], dotarray[57][98], dotarray[58][98], dotarray[59][98], dotarray[60][98], dotarray[61][98], dotarray[62][98], dotarray[63][98], dotarray[64][98], dotarray[65][98], dotarray[66][98], dotarray[67][98], dotarray[68][98], dotarray[69][98], dotarray[70][98], dotarray[71][98], dotarray[72][98], dotarray[73][98], dotarray[74][98], dotarray[75][98], dotarray[76][98], dotarray[77][98], dotarray[78][98], dotarray[79][98], dotarray[80][98], dotarray[81][98], dotarray[82][98], dotarray[83][98], dotarray[84][98], dotarray[85][98], dotarray[86][98], dotarray[87][98], dotarray[88][98], dotarray[89][98], dotarray[90][98], dotarray[91][98], dotarray[92][98], dotarray[93][98], dotarray[94][98], dotarray[95][98], dotarray[96][98], dotarray[97][98], dotarray[98][98], dotarray[99][98], dotarray[100][98], dotarray[101][98], dotarray[102][98], dotarray[103][98], dotarray[104][98], dotarray[105][98], dotarray[106][98], dotarray[107][98], dotarray[108][98], dotarray[109][98], dotarray[110][98], dotarray[111][98], dotarray[112][98], dotarray[113][98], dotarray[114][98], dotarray[115][98], dotarray[116][98], dotarray[117][98], dotarray[118][98], dotarray[119][98], dotarray[120][98], dotarray[121][98], dotarray[122][98], dotarray[123][98], dotarray[124][98], dotarray[125][98], dotarray[126][98], dotarray[127][98]};
assign dot_col_99 = {dotarray[0][99], dotarray[1][99], dotarray[2][99], dotarray[3][99], dotarray[4][99], dotarray[5][99], dotarray[6][99], dotarray[7][99], dotarray[8][99], dotarray[9][99], dotarray[10][99], dotarray[11][99], dotarray[12][99], dotarray[13][99], dotarray[14][99], dotarray[15][99], dotarray[16][99], dotarray[17][99], dotarray[18][99], dotarray[19][99], dotarray[20][99], dotarray[21][99], dotarray[22][99], dotarray[23][99], dotarray[24][99], dotarray[25][99], dotarray[26][99], dotarray[27][99], dotarray[28][99], dotarray[29][99], dotarray[30][99], dotarray[31][99], dotarray[32][99], dotarray[33][99], dotarray[34][99], dotarray[35][99], dotarray[36][99], dotarray[37][99], dotarray[38][99], dotarray[39][99], dotarray[40][99], dotarray[41][99], dotarray[42][99], dotarray[43][99], dotarray[44][99], dotarray[45][99], dotarray[46][99], dotarray[47][99], dotarray[48][99], dotarray[49][99], dotarray[50][99], dotarray[51][99], dotarray[52][99], dotarray[53][99], dotarray[54][99], dotarray[55][99], dotarray[56][99], dotarray[57][99], dotarray[58][99], dotarray[59][99], dotarray[60][99], dotarray[61][99], dotarray[62][99], dotarray[63][99], dotarray[64][99], dotarray[65][99], dotarray[66][99], dotarray[67][99], dotarray[68][99], dotarray[69][99], dotarray[70][99], dotarray[71][99], dotarray[72][99], dotarray[73][99], dotarray[74][99], dotarray[75][99], dotarray[76][99], dotarray[77][99], dotarray[78][99], dotarray[79][99], dotarray[80][99], dotarray[81][99], dotarray[82][99], dotarray[83][99], dotarray[84][99], dotarray[85][99], dotarray[86][99], dotarray[87][99], dotarray[88][99], dotarray[89][99], dotarray[90][99], dotarray[91][99], dotarray[92][99], dotarray[93][99], dotarray[94][99], dotarray[95][99], dotarray[96][99], dotarray[97][99], dotarray[98][99], dotarray[99][99], dotarray[100][99], dotarray[101][99], dotarray[102][99], dotarray[103][99], dotarray[104][99], dotarray[105][99], dotarray[106][99], dotarray[107][99], dotarray[108][99], dotarray[109][99], dotarray[110][99], dotarray[111][99], dotarray[112][99], dotarray[113][99], dotarray[114][99], dotarray[115][99], dotarray[116][99], dotarray[117][99], dotarray[118][99], dotarray[119][99], dotarray[120][99], dotarray[121][99], dotarray[122][99], dotarray[123][99], dotarray[124][99], dotarray[125][99], dotarray[126][99], dotarray[127][99]};
assign dot_col_100 = {dotarray[0][100], dotarray[1][100], dotarray[2][100], dotarray[3][100], dotarray[4][100], dotarray[5][100], dotarray[6][100], dotarray[7][100], dotarray[8][100], dotarray[9][100], dotarray[10][100], dotarray[11][100], dotarray[12][100], dotarray[13][100], dotarray[14][100], dotarray[15][100], dotarray[16][100], dotarray[17][100], dotarray[18][100], dotarray[19][100], dotarray[20][100], dotarray[21][100], dotarray[22][100], dotarray[23][100], dotarray[24][100], dotarray[25][100], dotarray[26][100], dotarray[27][100], dotarray[28][100], dotarray[29][100], dotarray[30][100], dotarray[31][100], dotarray[32][100], dotarray[33][100], dotarray[34][100], dotarray[35][100], dotarray[36][100], dotarray[37][100], dotarray[38][100], dotarray[39][100], dotarray[40][100], dotarray[41][100], dotarray[42][100], dotarray[43][100], dotarray[44][100], dotarray[45][100], dotarray[46][100], dotarray[47][100], dotarray[48][100], dotarray[49][100], dotarray[50][100], dotarray[51][100], dotarray[52][100], dotarray[53][100], dotarray[54][100], dotarray[55][100], dotarray[56][100], dotarray[57][100], dotarray[58][100], dotarray[59][100], dotarray[60][100], dotarray[61][100], dotarray[62][100], dotarray[63][100], dotarray[64][100], dotarray[65][100], dotarray[66][100], dotarray[67][100], dotarray[68][100], dotarray[69][100], dotarray[70][100], dotarray[71][100], dotarray[72][100], dotarray[73][100], dotarray[74][100], dotarray[75][100], dotarray[76][100], dotarray[77][100], dotarray[78][100], dotarray[79][100], dotarray[80][100], dotarray[81][100], dotarray[82][100], dotarray[83][100], dotarray[84][100], dotarray[85][100], dotarray[86][100], dotarray[87][100], dotarray[88][100], dotarray[89][100], dotarray[90][100], dotarray[91][100], dotarray[92][100], dotarray[93][100], dotarray[94][100], dotarray[95][100], dotarray[96][100], dotarray[97][100], dotarray[98][100], dotarray[99][100], dotarray[100][100], dotarray[101][100], dotarray[102][100], dotarray[103][100], dotarray[104][100], dotarray[105][100], dotarray[106][100], dotarray[107][100], dotarray[108][100], dotarray[109][100], dotarray[110][100], dotarray[111][100], dotarray[112][100], dotarray[113][100], dotarray[114][100], dotarray[115][100], dotarray[116][100], dotarray[117][100], dotarray[118][100], dotarray[119][100], dotarray[120][100], dotarray[121][100], dotarray[122][100], dotarray[123][100], dotarray[124][100], dotarray[125][100], dotarray[126][100], dotarray[127][100]};
assign dot_col_101 = {dotarray[0][101], dotarray[1][101], dotarray[2][101], dotarray[3][101], dotarray[4][101], dotarray[5][101], dotarray[6][101], dotarray[7][101], dotarray[8][101], dotarray[9][101], dotarray[10][101], dotarray[11][101], dotarray[12][101], dotarray[13][101], dotarray[14][101], dotarray[15][101], dotarray[16][101], dotarray[17][101], dotarray[18][101], dotarray[19][101], dotarray[20][101], dotarray[21][101], dotarray[22][101], dotarray[23][101], dotarray[24][101], dotarray[25][101], dotarray[26][101], dotarray[27][101], dotarray[28][101], dotarray[29][101], dotarray[30][101], dotarray[31][101], dotarray[32][101], dotarray[33][101], dotarray[34][101], dotarray[35][101], dotarray[36][101], dotarray[37][101], dotarray[38][101], dotarray[39][101], dotarray[40][101], dotarray[41][101], dotarray[42][101], dotarray[43][101], dotarray[44][101], dotarray[45][101], dotarray[46][101], dotarray[47][101], dotarray[48][101], dotarray[49][101], dotarray[50][101], dotarray[51][101], dotarray[52][101], dotarray[53][101], dotarray[54][101], dotarray[55][101], dotarray[56][101], dotarray[57][101], dotarray[58][101], dotarray[59][101], dotarray[60][101], dotarray[61][101], dotarray[62][101], dotarray[63][101], dotarray[64][101], dotarray[65][101], dotarray[66][101], dotarray[67][101], dotarray[68][101], dotarray[69][101], dotarray[70][101], dotarray[71][101], dotarray[72][101], dotarray[73][101], dotarray[74][101], dotarray[75][101], dotarray[76][101], dotarray[77][101], dotarray[78][101], dotarray[79][101], dotarray[80][101], dotarray[81][101], dotarray[82][101], dotarray[83][101], dotarray[84][101], dotarray[85][101], dotarray[86][101], dotarray[87][101], dotarray[88][101], dotarray[89][101], dotarray[90][101], dotarray[91][101], dotarray[92][101], dotarray[93][101], dotarray[94][101], dotarray[95][101], dotarray[96][101], dotarray[97][101], dotarray[98][101], dotarray[99][101], dotarray[100][101], dotarray[101][101], dotarray[102][101], dotarray[103][101], dotarray[104][101], dotarray[105][101], dotarray[106][101], dotarray[107][101], dotarray[108][101], dotarray[109][101], dotarray[110][101], dotarray[111][101], dotarray[112][101], dotarray[113][101], dotarray[114][101], dotarray[115][101], dotarray[116][101], dotarray[117][101], dotarray[118][101], dotarray[119][101], dotarray[120][101], dotarray[121][101], dotarray[122][101], dotarray[123][101], dotarray[124][101], dotarray[125][101], dotarray[126][101], dotarray[127][101]};
assign dot_col_102 = {dotarray[0][102], dotarray[1][102], dotarray[2][102], dotarray[3][102], dotarray[4][102], dotarray[5][102], dotarray[6][102], dotarray[7][102], dotarray[8][102], dotarray[9][102], dotarray[10][102], dotarray[11][102], dotarray[12][102], dotarray[13][102], dotarray[14][102], dotarray[15][102], dotarray[16][102], dotarray[17][102], dotarray[18][102], dotarray[19][102], dotarray[20][102], dotarray[21][102], dotarray[22][102], dotarray[23][102], dotarray[24][102], dotarray[25][102], dotarray[26][102], dotarray[27][102], dotarray[28][102], dotarray[29][102], dotarray[30][102], dotarray[31][102], dotarray[32][102], dotarray[33][102], dotarray[34][102], dotarray[35][102], dotarray[36][102], dotarray[37][102], dotarray[38][102], dotarray[39][102], dotarray[40][102], dotarray[41][102], dotarray[42][102], dotarray[43][102], dotarray[44][102], dotarray[45][102], dotarray[46][102], dotarray[47][102], dotarray[48][102], dotarray[49][102], dotarray[50][102], dotarray[51][102], dotarray[52][102], dotarray[53][102], dotarray[54][102], dotarray[55][102], dotarray[56][102], dotarray[57][102], dotarray[58][102], dotarray[59][102], dotarray[60][102], dotarray[61][102], dotarray[62][102], dotarray[63][102], dotarray[64][102], dotarray[65][102], dotarray[66][102], dotarray[67][102], dotarray[68][102], dotarray[69][102], dotarray[70][102], dotarray[71][102], dotarray[72][102], dotarray[73][102], dotarray[74][102], dotarray[75][102], dotarray[76][102], dotarray[77][102], dotarray[78][102], dotarray[79][102], dotarray[80][102], dotarray[81][102], dotarray[82][102], dotarray[83][102], dotarray[84][102], dotarray[85][102], dotarray[86][102], dotarray[87][102], dotarray[88][102], dotarray[89][102], dotarray[90][102], dotarray[91][102], dotarray[92][102], dotarray[93][102], dotarray[94][102], dotarray[95][102], dotarray[96][102], dotarray[97][102], dotarray[98][102], dotarray[99][102], dotarray[100][102], dotarray[101][102], dotarray[102][102], dotarray[103][102], dotarray[104][102], dotarray[105][102], dotarray[106][102], dotarray[107][102], dotarray[108][102], dotarray[109][102], dotarray[110][102], dotarray[111][102], dotarray[112][102], dotarray[113][102], dotarray[114][102], dotarray[115][102], dotarray[116][102], dotarray[117][102], dotarray[118][102], dotarray[119][102], dotarray[120][102], dotarray[121][102], dotarray[122][102], dotarray[123][102], dotarray[124][102], dotarray[125][102], dotarray[126][102], dotarray[127][102]};
assign dot_col_103 = {dotarray[0][103], dotarray[1][103], dotarray[2][103], dotarray[3][103], dotarray[4][103], dotarray[5][103], dotarray[6][103], dotarray[7][103], dotarray[8][103], dotarray[9][103], dotarray[10][103], dotarray[11][103], dotarray[12][103], dotarray[13][103], dotarray[14][103], dotarray[15][103], dotarray[16][103], dotarray[17][103], dotarray[18][103], dotarray[19][103], dotarray[20][103], dotarray[21][103], dotarray[22][103], dotarray[23][103], dotarray[24][103], dotarray[25][103], dotarray[26][103], dotarray[27][103], dotarray[28][103], dotarray[29][103], dotarray[30][103], dotarray[31][103], dotarray[32][103], dotarray[33][103], dotarray[34][103], dotarray[35][103], dotarray[36][103], dotarray[37][103], dotarray[38][103], dotarray[39][103], dotarray[40][103], dotarray[41][103], dotarray[42][103], dotarray[43][103], dotarray[44][103], dotarray[45][103], dotarray[46][103], dotarray[47][103], dotarray[48][103], dotarray[49][103], dotarray[50][103], dotarray[51][103], dotarray[52][103], dotarray[53][103], dotarray[54][103], dotarray[55][103], dotarray[56][103], dotarray[57][103], dotarray[58][103], dotarray[59][103], dotarray[60][103], dotarray[61][103], dotarray[62][103], dotarray[63][103], dotarray[64][103], dotarray[65][103], dotarray[66][103], dotarray[67][103], dotarray[68][103], dotarray[69][103], dotarray[70][103], dotarray[71][103], dotarray[72][103], dotarray[73][103], dotarray[74][103], dotarray[75][103], dotarray[76][103], dotarray[77][103], dotarray[78][103], dotarray[79][103], dotarray[80][103], dotarray[81][103], dotarray[82][103], dotarray[83][103], dotarray[84][103], dotarray[85][103], dotarray[86][103], dotarray[87][103], dotarray[88][103], dotarray[89][103], dotarray[90][103], dotarray[91][103], dotarray[92][103], dotarray[93][103], dotarray[94][103], dotarray[95][103], dotarray[96][103], dotarray[97][103], dotarray[98][103], dotarray[99][103], dotarray[100][103], dotarray[101][103], dotarray[102][103], dotarray[103][103], dotarray[104][103], dotarray[105][103], dotarray[106][103], dotarray[107][103], dotarray[108][103], dotarray[109][103], dotarray[110][103], dotarray[111][103], dotarray[112][103], dotarray[113][103], dotarray[114][103], dotarray[115][103], dotarray[116][103], dotarray[117][103], dotarray[118][103], dotarray[119][103], dotarray[120][103], dotarray[121][103], dotarray[122][103], dotarray[123][103], dotarray[124][103], dotarray[125][103], dotarray[126][103], dotarray[127][103]};
assign dot_col_104 = {dotarray[0][104], dotarray[1][104], dotarray[2][104], dotarray[3][104], dotarray[4][104], dotarray[5][104], dotarray[6][104], dotarray[7][104], dotarray[8][104], dotarray[9][104], dotarray[10][104], dotarray[11][104], dotarray[12][104], dotarray[13][104], dotarray[14][104], dotarray[15][104], dotarray[16][104], dotarray[17][104], dotarray[18][104], dotarray[19][104], dotarray[20][104], dotarray[21][104], dotarray[22][104], dotarray[23][104], dotarray[24][104], dotarray[25][104], dotarray[26][104], dotarray[27][104], dotarray[28][104], dotarray[29][104], dotarray[30][104], dotarray[31][104], dotarray[32][104], dotarray[33][104], dotarray[34][104], dotarray[35][104], dotarray[36][104], dotarray[37][104], dotarray[38][104], dotarray[39][104], dotarray[40][104], dotarray[41][104], dotarray[42][104], dotarray[43][104], dotarray[44][104], dotarray[45][104], dotarray[46][104], dotarray[47][104], dotarray[48][104], dotarray[49][104], dotarray[50][104], dotarray[51][104], dotarray[52][104], dotarray[53][104], dotarray[54][104], dotarray[55][104], dotarray[56][104], dotarray[57][104], dotarray[58][104], dotarray[59][104], dotarray[60][104], dotarray[61][104], dotarray[62][104], dotarray[63][104], dotarray[64][104], dotarray[65][104], dotarray[66][104], dotarray[67][104], dotarray[68][104], dotarray[69][104], dotarray[70][104], dotarray[71][104], dotarray[72][104], dotarray[73][104], dotarray[74][104], dotarray[75][104], dotarray[76][104], dotarray[77][104], dotarray[78][104], dotarray[79][104], dotarray[80][104], dotarray[81][104], dotarray[82][104], dotarray[83][104], dotarray[84][104], dotarray[85][104], dotarray[86][104], dotarray[87][104], dotarray[88][104], dotarray[89][104], dotarray[90][104], dotarray[91][104], dotarray[92][104], dotarray[93][104], dotarray[94][104], dotarray[95][104], dotarray[96][104], dotarray[97][104], dotarray[98][104], dotarray[99][104], dotarray[100][104], dotarray[101][104], dotarray[102][104], dotarray[103][104], dotarray[104][104], dotarray[105][104], dotarray[106][104], dotarray[107][104], dotarray[108][104], dotarray[109][104], dotarray[110][104], dotarray[111][104], dotarray[112][104], dotarray[113][104], dotarray[114][104], dotarray[115][104], dotarray[116][104], dotarray[117][104], dotarray[118][104], dotarray[119][104], dotarray[120][104], dotarray[121][104], dotarray[122][104], dotarray[123][104], dotarray[124][104], dotarray[125][104], dotarray[126][104], dotarray[127][104]};
assign dot_col_105 = {dotarray[0][105], dotarray[1][105], dotarray[2][105], dotarray[3][105], dotarray[4][105], dotarray[5][105], dotarray[6][105], dotarray[7][105], dotarray[8][105], dotarray[9][105], dotarray[10][105], dotarray[11][105], dotarray[12][105], dotarray[13][105], dotarray[14][105], dotarray[15][105], dotarray[16][105], dotarray[17][105], dotarray[18][105], dotarray[19][105], dotarray[20][105], dotarray[21][105], dotarray[22][105], dotarray[23][105], dotarray[24][105], dotarray[25][105], dotarray[26][105], dotarray[27][105], dotarray[28][105], dotarray[29][105], dotarray[30][105], dotarray[31][105], dotarray[32][105], dotarray[33][105], dotarray[34][105], dotarray[35][105], dotarray[36][105], dotarray[37][105], dotarray[38][105], dotarray[39][105], dotarray[40][105], dotarray[41][105], dotarray[42][105], dotarray[43][105], dotarray[44][105], dotarray[45][105], dotarray[46][105], dotarray[47][105], dotarray[48][105], dotarray[49][105], dotarray[50][105], dotarray[51][105], dotarray[52][105], dotarray[53][105], dotarray[54][105], dotarray[55][105], dotarray[56][105], dotarray[57][105], dotarray[58][105], dotarray[59][105], dotarray[60][105], dotarray[61][105], dotarray[62][105], dotarray[63][105], dotarray[64][105], dotarray[65][105], dotarray[66][105], dotarray[67][105], dotarray[68][105], dotarray[69][105], dotarray[70][105], dotarray[71][105], dotarray[72][105], dotarray[73][105], dotarray[74][105], dotarray[75][105], dotarray[76][105], dotarray[77][105], dotarray[78][105], dotarray[79][105], dotarray[80][105], dotarray[81][105], dotarray[82][105], dotarray[83][105], dotarray[84][105], dotarray[85][105], dotarray[86][105], dotarray[87][105], dotarray[88][105], dotarray[89][105], dotarray[90][105], dotarray[91][105], dotarray[92][105], dotarray[93][105], dotarray[94][105], dotarray[95][105], dotarray[96][105], dotarray[97][105], dotarray[98][105], dotarray[99][105], dotarray[100][105], dotarray[101][105], dotarray[102][105], dotarray[103][105], dotarray[104][105], dotarray[105][105], dotarray[106][105], dotarray[107][105], dotarray[108][105], dotarray[109][105], dotarray[110][105], dotarray[111][105], dotarray[112][105], dotarray[113][105], dotarray[114][105], dotarray[115][105], dotarray[116][105], dotarray[117][105], dotarray[118][105], dotarray[119][105], dotarray[120][105], dotarray[121][105], dotarray[122][105], dotarray[123][105], dotarray[124][105], dotarray[125][105], dotarray[126][105], dotarray[127][105]};
assign dot_col_106 = {dotarray[0][106], dotarray[1][106], dotarray[2][106], dotarray[3][106], dotarray[4][106], dotarray[5][106], dotarray[6][106], dotarray[7][106], dotarray[8][106], dotarray[9][106], dotarray[10][106], dotarray[11][106], dotarray[12][106], dotarray[13][106], dotarray[14][106], dotarray[15][106], dotarray[16][106], dotarray[17][106], dotarray[18][106], dotarray[19][106], dotarray[20][106], dotarray[21][106], dotarray[22][106], dotarray[23][106], dotarray[24][106], dotarray[25][106], dotarray[26][106], dotarray[27][106], dotarray[28][106], dotarray[29][106], dotarray[30][106], dotarray[31][106], dotarray[32][106], dotarray[33][106], dotarray[34][106], dotarray[35][106], dotarray[36][106], dotarray[37][106], dotarray[38][106], dotarray[39][106], dotarray[40][106], dotarray[41][106], dotarray[42][106], dotarray[43][106], dotarray[44][106], dotarray[45][106], dotarray[46][106], dotarray[47][106], dotarray[48][106], dotarray[49][106], dotarray[50][106], dotarray[51][106], dotarray[52][106], dotarray[53][106], dotarray[54][106], dotarray[55][106], dotarray[56][106], dotarray[57][106], dotarray[58][106], dotarray[59][106], dotarray[60][106], dotarray[61][106], dotarray[62][106], dotarray[63][106], dotarray[64][106], dotarray[65][106], dotarray[66][106], dotarray[67][106], dotarray[68][106], dotarray[69][106], dotarray[70][106], dotarray[71][106], dotarray[72][106], dotarray[73][106], dotarray[74][106], dotarray[75][106], dotarray[76][106], dotarray[77][106], dotarray[78][106], dotarray[79][106], dotarray[80][106], dotarray[81][106], dotarray[82][106], dotarray[83][106], dotarray[84][106], dotarray[85][106], dotarray[86][106], dotarray[87][106], dotarray[88][106], dotarray[89][106], dotarray[90][106], dotarray[91][106], dotarray[92][106], dotarray[93][106], dotarray[94][106], dotarray[95][106], dotarray[96][106], dotarray[97][106], dotarray[98][106], dotarray[99][106], dotarray[100][106], dotarray[101][106], dotarray[102][106], dotarray[103][106], dotarray[104][106], dotarray[105][106], dotarray[106][106], dotarray[107][106], dotarray[108][106], dotarray[109][106], dotarray[110][106], dotarray[111][106], dotarray[112][106], dotarray[113][106], dotarray[114][106], dotarray[115][106], dotarray[116][106], dotarray[117][106], dotarray[118][106], dotarray[119][106], dotarray[120][106], dotarray[121][106], dotarray[122][106], dotarray[123][106], dotarray[124][106], dotarray[125][106], dotarray[126][106], dotarray[127][106]};
assign dot_col_107 = {dotarray[0][107], dotarray[1][107], dotarray[2][107], dotarray[3][107], dotarray[4][107], dotarray[5][107], dotarray[6][107], dotarray[7][107], dotarray[8][107], dotarray[9][107], dotarray[10][107], dotarray[11][107], dotarray[12][107], dotarray[13][107], dotarray[14][107], dotarray[15][107], dotarray[16][107], dotarray[17][107], dotarray[18][107], dotarray[19][107], dotarray[20][107], dotarray[21][107], dotarray[22][107], dotarray[23][107], dotarray[24][107], dotarray[25][107], dotarray[26][107], dotarray[27][107], dotarray[28][107], dotarray[29][107], dotarray[30][107], dotarray[31][107], dotarray[32][107], dotarray[33][107], dotarray[34][107], dotarray[35][107], dotarray[36][107], dotarray[37][107], dotarray[38][107], dotarray[39][107], dotarray[40][107], dotarray[41][107], dotarray[42][107], dotarray[43][107], dotarray[44][107], dotarray[45][107], dotarray[46][107], dotarray[47][107], dotarray[48][107], dotarray[49][107], dotarray[50][107], dotarray[51][107], dotarray[52][107], dotarray[53][107], dotarray[54][107], dotarray[55][107], dotarray[56][107], dotarray[57][107], dotarray[58][107], dotarray[59][107], dotarray[60][107], dotarray[61][107], dotarray[62][107], dotarray[63][107], dotarray[64][107], dotarray[65][107], dotarray[66][107], dotarray[67][107], dotarray[68][107], dotarray[69][107], dotarray[70][107], dotarray[71][107], dotarray[72][107], dotarray[73][107], dotarray[74][107], dotarray[75][107], dotarray[76][107], dotarray[77][107], dotarray[78][107], dotarray[79][107], dotarray[80][107], dotarray[81][107], dotarray[82][107], dotarray[83][107], dotarray[84][107], dotarray[85][107], dotarray[86][107], dotarray[87][107], dotarray[88][107], dotarray[89][107], dotarray[90][107], dotarray[91][107], dotarray[92][107], dotarray[93][107], dotarray[94][107], dotarray[95][107], dotarray[96][107], dotarray[97][107], dotarray[98][107], dotarray[99][107], dotarray[100][107], dotarray[101][107], dotarray[102][107], dotarray[103][107], dotarray[104][107], dotarray[105][107], dotarray[106][107], dotarray[107][107], dotarray[108][107], dotarray[109][107], dotarray[110][107], dotarray[111][107], dotarray[112][107], dotarray[113][107], dotarray[114][107], dotarray[115][107], dotarray[116][107], dotarray[117][107], dotarray[118][107], dotarray[119][107], dotarray[120][107], dotarray[121][107], dotarray[122][107], dotarray[123][107], dotarray[124][107], dotarray[125][107], dotarray[126][107], dotarray[127][107]};
assign dot_col_108 = {dotarray[0][108], dotarray[1][108], dotarray[2][108], dotarray[3][108], dotarray[4][108], dotarray[5][108], dotarray[6][108], dotarray[7][108], dotarray[8][108], dotarray[9][108], dotarray[10][108], dotarray[11][108], dotarray[12][108], dotarray[13][108], dotarray[14][108], dotarray[15][108], dotarray[16][108], dotarray[17][108], dotarray[18][108], dotarray[19][108], dotarray[20][108], dotarray[21][108], dotarray[22][108], dotarray[23][108], dotarray[24][108], dotarray[25][108], dotarray[26][108], dotarray[27][108], dotarray[28][108], dotarray[29][108], dotarray[30][108], dotarray[31][108], dotarray[32][108], dotarray[33][108], dotarray[34][108], dotarray[35][108], dotarray[36][108], dotarray[37][108], dotarray[38][108], dotarray[39][108], dotarray[40][108], dotarray[41][108], dotarray[42][108], dotarray[43][108], dotarray[44][108], dotarray[45][108], dotarray[46][108], dotarray[47][108], dotarray[48][108], dotarray[49][108], dotarray[50][108], dotarray[51][108], dotarray[52][108], dotarray[53][108], dotarray[54][108], dotarray[55][108], dotarray[56][108], dotarray[57][108], dotarray[58][108], dotarray[59][108], dotarray[60][108], dotarray[61][108], dotarray[62][108], dotarray[63][108], dotarray[64][108], dotarray[65][108], dotarray[66][108], dotarray[67][108], dotarray[68][108], dotarray[69][108], dotarray[70][108], dotarray[71][108], dotarray[72][108], dotarray[73][108], dotarray[74][108], dotarray[75][108], dotarray[76][108], dotarray[77][108], dotarray[78][108], dotarray[79][108], dotarray[80][108], dotarray[81][108], dotarray[82][108], dotarray[83][108], dotarray[84][108], dotarray[85][108], dotarray[86][108], dotarray[87][108], dotarray[88][108], dotarray[89][108], dotarray[90][108], dotarray[91][108], dotarray[92][108], dotarray[93][108], dotarray[94][108], dotarray[95][108], dotarray[96][108], dotarray[97][108], dotarray[98][108], dotarray[99][108], dotarray[100][108], dotarray[101][108], dotarray[102][108], dotarray[103][108], dotarray[104][108], dotarray[105][108], dotarray[106][108], dotarray[107][108], dotarray[108][108], dotarray[109][108], dotarray[110][108], dotarray[111][108], dotarray[112][108], dotarray[113][108], dotarray[114][108], dotarray[115][108], dotarray[116][108], dotarray[117][108], dotarray[118][108], dotarray[119][108], dotarray[120][108], dotarray[121][108], dotarray[122][108], dotarray[123][108], dotarray[124][108], dotarray[125][108], dotarray[126][108], dotarray[127][108]};
assign dot_col_109 = {dotarray[0][109], dotarray[1][109], dotarray[2][109], dotarray[3][109], dotarray[4][109], dotarray[5][109], dotarray[6][109], dotarray[7][109], dotarray[8][109], dotarray[9][109], dotarray[10][109], dotarray[11][109], dotarray[12][109], dotarray[13][109], dotarray[14][109], dotarray[15][109], dotarray[16][109], dotarray[17][109], dotarray[18][109], dotarray[19][109], dotarray[20][109], dotarray[21][109], dotarray[22][109], dotarray[23][109], dotarray[24][109], dotarray[25][109], dotarray[26][109], dotarray[27][109], dotarray[28][109], dotarray[29][109], dotarray[30][109], dotarray[31][109], dotarray[32][109], dotarray[33][109], dotarray[34][109], dotarray[35][109], dotarray[36][109], dotarray[37][109], dotarray[38][109], dotarray[39][109], dotarray[40][109], dotarray[41][109], dotarray[42][109], dotarray[43][109], dotarray[44][109], dotarray[45][109], dotarray[46][109], dotarray[47][109], dotarray[48][109], dotarray[49][109], dotarray[50][109], dotarray[51][109], dotarray[52][109], dotarray[53][109], dotarray[54][109], dotarray[55][109], dotarray[56][109], dotarray[57][109], dotarray[58][109], dotarray[59][109], dotarray[60][109], dotarray[61][109], dotarray[62][109], dotarray[63][109], dotarray[64][109], dotarray[65][109], dotarray[66][109], dotarray[67][109], dotarray[68][109], dotarray[69][109], dotarray[70][109], dotarray[71][109], dotarray[72][109], dotarray[73][109], dotarray[74][109], dotarray[75][109], dotarray[76][109], dotarray[77][109], dotarray[78][109], dotarray[79][109], dotarray[80][109], dotarray[81][109], dotarray[82][109], dotarray[83][109], dotarray[84][109], dotarray[85][109], dotarray[86][109], dotarray[87][109], dotarray[88][109], dotarray[89][109], dotarray[90][109], dotarray[91][109], dotarray[92][109], dotarray[93][109], dotarray[94][109], dotarray[95][109], dotarray[96][109], dotarray[97][109], dotarray[98][109], dotarray[99][109], dotarray[100][109], dotarray[101][109], dotarray[102][109], dotarray[103][109], dotarray[104][109], dotarray[105][109], dotarray[106][109], dotarray[107][109], dotarray[108][109], dotarray[109][109], dotarray[110][109], dotarray[111][109], dotarray[112][109], dotarray[113][109], dotarray[114][109], dotarray[115][109], dotarray[116][109], dotarray[117][109], dotarray[118][109], dotarray[119][109], dotarray[120][109], dotarray[121][109], dotarray[122][109], dotarray[123][109], dotarray[124][109], dotarray[125][109], dotarray[126][109], dotarray[127][109]};
assign dot_col_110 = {dotarray[0][110], dotarray[1][110], dotarray[2][110], dotarray[3][110], dotarray[4][110], dotarray[5][110], dotarray[6][110], dotarray[7][110], dotarray[8][110], dotarray[9][110], dotarray[10][110], dotarray[11][110], dotarray[12][110], dotarray[13][110], dotarray[14][110], dotarray[15][110], dotarray[16][110], dotarray[17][110], dotarray[18][110], dotarray[19][110], dotarray[20][110], dotarray[21][110], dotarray[22][110], dotarray[23][110], dotarray[24][110], dotarray[25][110], dotarray[26][110], dotarray[27][110], dotarray[28][110], dotarray[29][110], dotarray[30][110], dotarray[31][110], dotarray[32][110], dotarray[33][110], dotarray[34][110], dotarray[35][110], dotarray[36][110], dotarray[37][110], dotarray[38][110], dotarray[39][110], dotarray[40][110], dotarray[41][110], dotarray[42][110], dotarray[43][110], dotarray[44][110], dotarray[45][110], dotarray[46][110], dotarray[47][110], dotarray[48][110], dotarray[49][110], dotarray[50][110], dotarray[51][110], dotarray[52][110], dotarray[53][110], dotarray[54][110], dotarray[55][110], dotarray[56][110], dotarray[57][110], dotarray[58][110], dotarray[59][110], dotarray[60][110], dotarray[61][110], dotarray[62][110], dotarray[63][110], dotarray[64][110], dotarray[65][110], dotarray[66][110], dotarray[67][110], dotarray[68][110], dotarray[69][110], dotarray[70][110], dotarray[71][110], dotarray[72][110], dotarray[73][110], dotarray[74][110], dotarray[75][110], dotarray[76][110], dotarray[77][110], dotarray[78][110], dotarray[79][110], dotarray[80][110], dotarray[81][110], dotarray[82][110], dotarray[83][110], dotarray[84][110], dotarray[85][110], dotarray[86][110], dotarray[87][110], dotarray[88][110], dotarray[89][110], dotarray[90][110], dotarray[91][110], dotarray[92][110], dotarray[93][110], dotarray[94][110], dotarray[95][110], dotarray[96][110], dotarray[97][110], dotarray[98][110], dotarray[99][110], dotarray[100][110], dotarray[101][110], dotarray[102][110], dotarray[103][110], dotarray[104][110], dotarray[105][110], dotarray[106][110], dotarray[107][110], dotarray[108][110], dotarray[109][110], dotarray[110][110], dotarray[111][110], dotarray[112][110], dotarray[113][110], dotarray[114][110], dotarray[115][110], dotarray[116][110], dotarray[117][110], dotarray[118][110], dotarray[119][110], dotarray[120][110], dotarray[121][110], dotarray[122][110], dotarray[123][110], dotarray[124][110], dotarray[125][110], dotarray[126][110], dotarray[127][110]};
assign dot_col_111 = {dotarray[0][111], dotarray[1][111], dotarray[2][111], dotarray[3][111], dotarray[4][111], dotarray[5][111], dotarray[6][111], dotarray[7][111], dotarray[8][111], dotarray[9][111], dotarray[10][111], dotarray[11][111], dotarray[12][111], dotarray[13][111], dotarray[14][111], dotarray[15][111], dotarray[16][111], dotarray[17][111], dotarray[18][111], dotarray[19][111], dotarray[20][111], dotarray[21][111], dotarray[22][111], dotarray[23][111], dotarray[24][111], dotarray[25][111], dotarray[26][111], dotarray[27][111], dotarray[28][111], dotarray[29][111], dotarray[30][111], dotarray[31][111], dotarray[32][111], dotarray[33][111], dotarray[34][111], dotarray[35][111], dotarray[36][111], dotarray[37][111], dotarray[38][111], dotarray[39][111], dotarray[40][111], dotarray[41][111], dotarray[42][111], dotarray[43][111], dotarray[44][111], dotarray[45][111], dotarray[46][111], dotarray[47][111], dotarray[48][111], dotarray[49][111], dotarray[50][111], dotarray[51][111], dotarray[52][111], dotarray[53][111], dotarray[54][111], dotarray[55][111], dotarray[56][111], dotarray[57][111], dotarray[58][111], dotarray[59][111], dotarray[60][111], dotarray[61][111], dotarray[62][111], dotarray[63][111], dotarray[64][111], dotarray[65][111], dotarray[66][111], dotarray[67][111], dotarray[68][111], dotarray[69][111], dotarray[70][111], dotarray[71][111], dotarray[72][111], dotarray[73][111], dotarray[74][111], dotarray[75][111], dotarray[76][111], dotarray[77][111], dotarray[78][111], dotarray[79][111], dotarray[80][111], dotarray[81][111], dotarray[82][111], dotarray[83][111], dotarray[84][111], dotarray[85][111], dotarray[86][111], dotarray[87][111], dotarray[88][111], dotarray[89][111], dotarray[90][111], dotarray[91][111], dotarray[92][111], dotarray[93][111], dotarray[94][111], dotarray[95][111], dotarray[96][111], dotarray[97][111], dotarray[98][111], dotarray[99][111], dotarray[100][111], dotarray[101][111], dotarray[102][111], dotarray[103][111], dotarray[104][111], dotarray[105][111], dotarray[106][111], dotarray[107][111], dotarray[108][111], dotarray[109][111], dotarray[110][111], dotarray[111][111], dotarray[112][111], dotarray[113][111], dotarray[114][111], dotarray[115][111], dotarray[116][111], dotarray[117][111], dotarray[118][111], dotarray[119][111], dotarray[120][111], dotarray[121][111], dotarray[122][111], dotarray[123][111], dotarray[124][111], dotarray[125][111], dotarray[126][111], dotarray[127][111]};
assign dot_col_112 = {dotarray[0][112], dotarray[1][112], dotarray[2][112], dotarray[3][112], dotarray[4][112], dotarray[5][112], dotarray[6][112], dotarray[7][112], dotarray[8][112], dotarray[9][112], dotarray[10][112], dotarray[11][112], dotarray[12][112], dotarray[13][112], dotarray[14][112], dotarray[15][112], dotarray[16][112], dotarray[17][112], dotarray[18][112], dotarray[19][112], dotarray[20][112], dotarray[21][112], dotarray[22][112], dotarray[23][112], dotarray[24][112], dotarray[25][112], dotarray[26][112], dotarray[27][112], dotarray[28][112], dotarray[29][112], dotarray[30][112], dotarray[31][112], dotarray[32][112], dotarray[33][112], dotarray[34][112], dotarray[35][112], dotarray[36][112], dotarray[37][112], dotarray[38][112], dotarray[39][112], dotarray[40][112], dotarray[41][112], dotarray[42][112], dotarray[43][112], dotarray[44][112], dotarray[45][112], dotarray[46][112], dotarray[47][112], dotarray[48][112], dotarray[49][112], dotarray[50][112], dotarray[51][112], dotarray[52][112], dotarray[53][112], dotarray[54][112], dotarray[55][112], dotarray[56][112], dotarray[57][112], dotarray[58][112], dotarray[59][112], dotarray[60][112], dotarray[61][112], dotarray[62][112], dotarray[63][112], dotarray[64][112], dotarray[65][112], dotarray[66][112], dotarray[67][112], dotarray[68][112], dotarray[69][112], dotarray[70][112], dotarray[71][112], dotarray[72][112], dotarray[73][112], dotarray[74][112], dotarray[75][112], dotarray[76][112], dotarray[77][112], dotarray[78][112], dotarray[79][112], dotarray[80][112], dotarray[81][112], dotarray[82][112], dotarray[83][112], dotarray[84][112], dotarray[85][112], dotarray[86][112], dotarray[87][112], dotarray[88][112], dotarray[89][112], dotarray[90][112], dotarray[91][112], dotarray[92][112], dotarray[93][112], dotarray[94][112], dotarray[95][112], dotarray[96][112], dotarray[97][112], dotarray[98][112], dotarray[99][112], dotarray[100][112], dotarray[101][112], dotarray[102][112], dotarray[103][112], dotarray[104][112], dotarray[105][112], dotarray[106][112], dotarray[107][112], dotarray[108][112], dotarray[109][112], dotarray[110][112], dotarray[111][112], dotarray[112][112], dotarray[113][112], dotarray[114][112], dotarray[115][112], dotarray[116][112], dotarray[117][112], dotarray[118][112], dotarray[119][112], dotarray[120][112], dotarray[121][112], dotarray[122][112], dotarray[123][112], dotarray[124][112], dotarray[125][112], dotarray[126][112], dotarray[127][112]};
assign dot_col_113 = {dotarray[0][113], dotarray[1][113], dotarray[2][113], dotarray[3][113], dotarray[4][113], dotarray[5][113], dotarray[6][113], dotarray[7][113], dotarray[8][113], dotarray[9][113], dotarray[10][113], dotarray[11][113], dotarray[12][113], dotarray[13][113], dotarray[14][113], dotarray[15][113], dotarray[16][113], dotarray[17][113], dotarray[18][113], dotarray[19][113], dotarray[20][113], dotarray[21][113], dotarray[22][113], dotarray[23][113], dotarray[24][113], dotarray[25][113], dotarray[26][113], dotarray[27][113], dotarray[28][113], dotarray[29][113], dotarray[30][113], dotarray[31][113], dotarray[32][113], dotarray[33][113], dotarray[34][113], dotarray[35][113], dotarray[36][113], dotarray[37][113], dotarray[38][113], dotarray[39][113], dotarray[40][113], dotarray[41][113], dotarray[42][113], dotarray[43][113], dotarray[44][113], dotarray[45][113], dotarray[46][113], dotarray[47][113], dotarray[48][113], dotarray[49][113], dotarray[50][113], dotarray[51][113], dotarray[52][113], dotarray[53][113], dotarray[54][113], dotarray[55][113], dotarray[56][113], dotarray[57][113], dotarray[58][113], dotarray[59][113], dotarray[60][113], dotarray[61][113], dotarray[62][113], dotarray[63][113], dotarray[64][113], dotarray[65][113], dotarray[66][113], dotarray[67][113], dotarray[68][113], dotarray[69][113], dotarray[70][113], dotarray[71][113], dotarray[72][113], dotarray[73][113], dotarray[74][113], dotarray[75][113], dotarray[76][113], dotarray[77][113], dotarray[78][113], dotarray[79][113], dotarray[80][113], dotarray[81][113], dotarray[82][113], dotarray[83][113], dotarray[84][113], dotarray[85][113], dotarray[86][113], dotarray[87][113], dotarray[88][113], dotarray[89][113], dotarray[90][113], dotarray[91][113], dotarray[92][113], dotarray[93][113], dotarray[94][113], dotarray[95][113], dotarray[96][113], dotarray[97][113], dotarray[98][113], dotarray[99][113], dotarray[100][113], dotarray[101][113], dotarray[102][113], dotarray[103][113], dotarray[104][113], dotarray[105][113], dotarray[106][113], dotarray[107][113], dotarray[108][113], dotarray[109][113], dotarray[110][113], dotarray[111][113], dotarray[112][113], dotarray[113][113], dotarray[114][113], dotarray[115][113], dotarray[116][113], dotarray[117][113], dotarray[118][113], dotarray[119][113], dotarray[120][113], dotarray[121][113], dotarray[122][113], dotarray[123][113], dotarray[124][113], dotarray[125][113], dotarray[126][113], dotarray[127][113]};
assign dot_col_114 = {dotarray[0][114], dotarray[1][114], dotarray[2][114], dotarray[3][114], dotarray[4][114], dotarray[5][114], dotarray[6][114], dotarray[7][114], dotarray[8][114], dotarray[9][114], dotarray[10][114], dotarray[11][114], dotarray[12][114], dotarray[13][114], dotarray[14][114], dotarray[15][114], dotarray[16][114], dotarray[17][114], dotarray[18][114], dotarray[19][114], dotarray[20][114], dotarray[21][114], dotarray[22][114], dotarray[23][114], dotarray[24][114], dotarray[25][114], dotarray[26][114], dotarray[27][114], dotarray[28][114], dotarray[29][114], dotarray[30][114], dotarray[31][114], dotarray[32][114], dotarray[33][114], dotarray[34][114], dotarray[35][114], dotarray[36][114], dotarray[37][114], dotarray[38][114], dotarray[39][114], dotarray[40][114], dotarray[41][114], dotarray[42][114], dotarray[43][114], dotarray[44][114], dotarray[45][114], dotarray[46][114], dotarray[47][114], dotarray[48][114], dotarray[49][114], dotarray[50][114], dotarray[51][114], dotarray[52][114], dotarray[53][114], dotarray[54][114], dotarray[55][114], dotarray[56][114], dotarray[57][114], dotarray[58][114], dotarray[59][114], dotarray[60][114], dotarray[61][114], dotarray[62][114], dotarray[63][114], dotarray[64][114], dotarray[65][114], dotarray[66][114], dotarray[67][114], dotarray[68][114], dotarray[69][114], dotarray[70][114], dotarray[71][114], dotarray[72][114], dotarray[73][114], dotarray[74][114], dotarray[75][114], dotarray[76][114], dotarray[77][114], dotarray[78][114], dotarray[79][114], dotarray[80][114], dotarray[81][114], dotarray[82][114], dotarray[83][114], dotarray[84][114], dotarray[85][114], dotarray[86][114], dotarray[87][114], dotarray[88][114], dotarray[89][114], dotarray[90][114], dotarray[91][114], dotarray[92][114], dotarray[93][114], dotarray[94][114], dotarray[95][114], dotarray[96][114], dotarray[97][114], dotarray[98][114], dotarray[99][114], dotarray[100][114], dotarray[101][114], dotarray[102][114], dotarray[103][114], dotarray[104][114], dotarray[105][114], dotarray[106][114], dotarray[107][114], dotarray[108][114], dotarray[109][114], dotarray[110][114], dotarray[111][114], dotarray[112][114], dotarray[113][114], dotarray[114][114], dotarray[115][114], dotarray[116][114], dotarray[117][114], dotarray[118][114], dotarray[119][114], dotarray[120][114], dotarray[121][114], dotarray[122][114], dotarray[123][114], dotarray[124][114], dotarray[125][114], dotarray[126][114], dotarray[127][114]};
assign dot_col_115 = {dotarray[0][115], dotarray[1][115], dotarray[2][115], dotarray[3][115], dotarray[4][115], dotarray[5][115], dotarray[6][115], dotarray[7][115], dotarray[8][115], dotarray[9][115], dotarray[10][115], dotarray[11][115], dotarray[12][115], dotarray[13][115], dotarray[14][115], dotarray[15][115], dotarray[16][115], dotarray[17][115], dotarray[18][115], dotarray[19][115], dotarray[20][115], dotarray[21][115], dotarray[22][115], dotarray[23][115], dotarray[24][115], dotarray[25][115], dotarray[26][115], dotarray[27][115], dotarray[28][115], dotarray[29][115], dotarray[30][115], dotarray[31][115], dotarray[32][115], dotarray[33][115], dotarray[34][115], dotarray[35][115], dotarray[36][115], dotarray[37][115], dotarray[38][115], dotarray[39][115], dotarray[40][115], dotarray[41][115], dotarray[42][115], dotarray[43][115], dotarray[44][115], dotarray[45][115], dotarray[46][115], dotarray[47][115], dotarray[48][115], dotarray[49][115], dotarray[50][115], dotarray[51][115], dotarray[52][115], dotarray[53][115], dotarray[54][115], dotarray[55][115], dotarray[56][115], dotarray[57][115], dotarray[58][115], dotarray[59][115], dotarray[60][115], dotarray[61][115], dotarray[62][115], dotarray[63][115], dotarray[64][115], dotarray[65][115], dotarray[66][115], dotarray[67][115], dotarray[68][115], dotarray[69][115], dotarray[70][115], dotarray[71][115], dotarray[72][115], dotarray[73][115], dotarray[74][115], dotarray[75][115], dotarray[76][115], dotarray[77][115], dotarray[78][115], dotarray[79][115], dotarray[80][115], dotarray[81][115], dotarray[82][115], dotarray[83][115], dotarray[84][115], dotarray[85][115], dotarray[86][115], dotarray[87][115], dotarray[88][115], dotarray[89][115], dotarray[90][115], dotarray[91][115], dotarray[92][115], dotarray[93][115], dotarray[94][115], dotarray[95][115], dotarray[96][115], dotarray[97][115], dotarray[98][115], dotarray[99][115], dotarray[100][115], dotarray[101][115], dotarray[102][115], dotarray[103][115], dotarray[104][115], dotarray[105][115], dotarray[106][115], dotarray[107][115], dotarray[108][115], dotarray[109][115], dotarray[110][115], dotarray[111][115], dotarray[112][115], dotarray[113][115], dotarray[114][115], dotarray[115][115], dotarray[116][115], dotarray[117][115], dotarray[118][115], dotarray[119][115], dotarray[120][115], dotarray[121][115], dotarray[122][115], dotarray[123][115], dotarray[124][115], dotarray[125][115], dotarray[126][115], dotarray[127][115]};
assign dot_col_116 = {dotarray[0][116], dotarray[1][116], dotarray[2][116], dotarray[3][116], dotarray[4][116], dotarray[5][116], dotarray[6][116], dotarray[7][116], dotarray[8][116], dotarray[9][116], dotarray[10][116], dotarray[11][116], dotarray[12][116], dotarray[13][116], dotarray[14][116], dotarray[15][116], dotarray[16][116], dotarray[17][116], dotarray[18][116], dotarray[19][116], dotarray[20][116], dotarray[21][116], dotarray[22][116], dotarray[23][116], dotarray[24][116], dotarray[25][116], dotarray[26][116], dotarray[27][116], dotarray[28][116], dotarray[29][116], dotarray[30][116], dotarray[31][116], dotarray[32][116], dotarray[33][116], dotarray[34][116], dotarray[35][116], dotarray[36][116], dotarray[37][116], dotarray[38][116], dotarray[39][116], dotarray[40][116], dotarray[41][116], dotarray[42][116], dotarray[43][116], dotarray[44][116], dotarray[45][116], dotarray[46][116], dotarray[47][116], dotarray[48][116], dotarray[49][116], dotarray[50][116], dotarray[51][116], dotarray[52][116], dotarray[53][116], dotarray[54][116], dotarray[55][116], dotarray[56][116], dotarray[57][116], dotarray[58][116], dotarray[59][116], dotarray[60][116], dotarray[61][116], dotarray[62][116], dotarray[63][116], dotarray[64][116], dotarray[65][116], dotarray[66][116], dotarray[67][116], dotarray[68][116], dotarray[69][116], dotarray[70][116], dotarray[71][116], dotarray[72][116], dotarray[73][116], dotarray[74][116], dotarray[75][116], dotarray[76][116], dotarray[77][116], dotarray[78][116], dotarray[79][116], dotarray[80][116], dotarray[81][116], dotarray[82][116], dotarray[83][116], dotarray[84][116], dotarray[85][116], dotarray[86][116], dotarray[87][116], dotarray[88][116], dotarray[89][116], dotarray[90][116], dotarray[91][116], dotarray[92][116], dotarray[93][116], dotarray[94][116], dotarray[95][116], dotarray[96][116], dotarray[97][116], dotarray[98][116], dotarray[99][116], dotarray[100][116], dotarray[101][116], dotarray[102][116], dotarray[103][116], dotarray[104][116], dotarray[105][116], dotarray[106][116], dotarray[107][116], dotarray[108][116], dotarray[109][116], dotarray[110][116], dotarray[111][116], dotarray[112][116], dotarray[113][116], dotarray[114][116], dotarray[115][116], dotarray[116][116], dotarray[117][116], dotarray[118][116], dotarray[119][116], dotarray[120][116], dotarray[121][116], dotarray[122][116], dotarray[123][116], dotarray[124][116], dotarray[125][116], dotarray[126][116], dotarray[127][116]};
assign dot_col_117 = {dotarray[0][117], dotarray[1][117], dotarray[2][117], dotarray[3][117], dotarray[4][117], dotarray[5][117], dotarray[6][117], dotarray[7][117], dotarray[8][117], dotarray[9][117], dotarray[10][117], dotarray[11][117], dotarray[12][117], dotarray[13][117], dotarray[14][117], dotarray[15][117], dotarray[16][117], dotarray[17][117], dotarray[18][117], dotarray[19][117], dotarray[20][117], dotarray[21][117], dotarray[22][117], dotarray[23][117], dotarray[24][117], dotarray[25][117], dotarray[26][117], dotarray[27][117], dotarray[28][117], dotarray[29][117], dotarray[30][117], dotarray[31][117], dotarray[32][117], dotarray[33][117], dotarray[34][117], dotarray[35][117], dotarray[36][117], dotarray[37][117], dotarray[38][117], dotarray[39][117], dotarray[40][117], dotarray[41][117], dotarray[42][117], dotarray[43][117], dotarray[44][117], dotarray[45][117], dotarray[46][117], dotarray[47][117], dotarray[48][117], dotarray[49][117], dotarray[50][117], dotarray[51][117], dotarray[52][117], dotarray[53][117], dotarray[54][117], dotarray[55][117], dotarray[56][117], dotarray[57][117], dotarray[58][117], dotarray[59][117], dotarray[60][117], dotarray[61][117], dotarray[62][117], dotarray[63][117], dotarray[64][117], dotarray[65][117], dotarray[66][117], dotarray[67][117], dotarray[68][117], dotarray[69][117], dotarray[70][117], dotarray[71][117], dotarray[72][117], dotarray[73][117], dotarray[74][117], dotarray[75][117], dotarray[76][117], dotarray[77][117], dotarray[78][117], dotarray[79][117], dotarray[80][117], dotarray[81][117], dotarray[82][117], dotarray[83][117], dotarray[84][117], dotarray[85][117], dotarray[86][117], dotarray[87][117], dotarray[88][117], dotarray[89][117], dotarray[90][117], dotarray[91][117], dotarray[92][117], dotarray[93][117], dotarray[94][117], dotarray[95][117], dotarray[96][117], dotarray[97][117], dotarray[98][117], dotarray[99][117], dotarray[100][117], dotarray[101][117], dotarray[102][117], dotarray[103][117], dotarray[104][117], dotarray[105][117], dotarray[106][117], dotarray[107][117], dotarray[108][117], dotarray[109][117], dotarray[110][117], dotarray[111][117], dotarray[112][117], dotarray[113][117], dotarray[114][117], dotarray[115][117], dotarray[116][117], dotarray[117][117], dotarray[118][117], dotarray[119][117], dotarray[120][117], dotarray[121][117], dotarray[122][117], dotarray[123][117], dotarray[124][117], dotarray[125][117], dotarray[126][117], dotarray[127][117]};
assign dot_col_118 = {dotarray[0][118], dotarray[1][118], dotarray[2][118], dotarray[3][118], dotarray[4][118], dotarray[5][118], dotarray[6][118], dotarray[7][118], dotarray[8][118], dotarray[9][118], dotarray[10][118], dotarray[11][118], dotarray[12][118], dotarray[13][118], dotarray[14][118], dotarray[15][118], dotarray[16][118], dotarray[17][118], dotarray[18][118], dotarray[19][118], dotarray[20][118], dotarray[21][118], dotarray[22][118], dotarray[23][118], dotarray[24][118], dotarray[25][118], dotarray[26][118], dotarray[27][118], dotarray[28][118], dotarray[29][118], dotarray[30][118], dotarray[31][118], dotarray[32][118], dotarray[33][118], dotarray[34][118], dotarray[35][118], dotarray[36][118], dotarray[37][118], dotarray[38][118], dotarray[39][118], dotarray[40][118], dotarray[41][118], dotarray[42][118], dotarray[43][118], dotarray[44][118], dotarray[45][118], dotarray[46][118], dotarray[47][118], dotarray[48][118], dotarray[49][118], dotarray[50][118], dotarray[51][118], dotarray[52][118], dotarray[53][118], dotarray[54][118], dotarray[55][118], dotarray[56][118], dotarray[57][118], dotarray[58][118], dotarray[59][118], dotarray[60][118], dotarray[61][118], dotarray[62][118], dotarray[63][118], dotarray[64][118], dotarray[65][118], dotarray[66][118], dotarray[67][118], dotarray[68][118], dotarray[69][118], dotarray[70][118], dotarray[71][118], dotarray[72][118], dotarray[73][118], dotarray[74][118], dotarray[75][118], dotarray[76][118], dotarray[77][118], dotarray[78][118], dotarray[79][118], dotarray[80][118], dotarray[81][118], dotarray[82][118], dotarray[83][118], dotarray[84][118], dotarray[85][118], dotarray[86][118], dotarray[87][118], dotarray[88][118], dotarray[89][118], dotarray[90][118], dotarray[91][118], dotarray[92][118], dotarray[93][118], dotarray[94][118], dotarray[95][118], dotarray[96][118], dotarray[97][118], dotarray[98][118], dotarray[99][118], dotarray[100][118], dotarray[101][118], dotarray[102][118], dotarray[103][118], dotarray[104][118], dotarray[105][118], dotarray[106][118], dotarray[107][118], dotarray[108][118], dotarray[109][118], dotarray[110][118], dotarray[111][118], dotarray[112][118], dotarray[113][118], dotarray[114][118], dotarray[115][118], dotarray[116][118], dotarray[117][118], dotarray[118][118], dotarray[119][118], dotarray[120][118], dotarray[121][118], dotarray[122][118], dotarray[123][118], dotarray[124][118], dotarray[125][118], dotarray[126][118], dotarray[127][118]};
assign dot_col_119 = {dotarray[0][119], dotarray[1][119], dotarray[2][119], dotarray[3][119], dotarray[4][119], dotarray[5][119], dotarray[6][119], dotarray[7][119], dotarray[8][119], dotarray[9][119], dotarray[10][119], dotarray[11][119], dotarray[12][119], dotarray[13][119], dotarray[14][119], dotarray[15][119], dotarray[16][119], dotarray[17][119], dotarray[18][119], dotarray[19][119], dotarray[20][119], dotarray[21][119], dotarray[22][119], dotarray[23][119], dotarray[24][119], dotarray[25][119], dotarray[26][119], dotarray[27][119], dotarray[28][119], dotarray[29][119], dotarray[30][119], dotarray[31][119], dotarray[32][119], dotarray[33][119], dotarray[34][119], dotarray[35][119], dotarray[36][119], dotarray[37][119], dotarray[38][119], dotarray[39][119], dotarray[40][119], dotarray[41][119], dotarray[42][119], dotarray[43][119], dotarray[44][119], dotarray[45][119], dotarray[46][119], dotarray[47][119], dotarray[48][119], dotarray[49][119], dotarray[50][119], dotarray[51][119], dotarray[52][119], dotarray[53][119], dotarray[54][119], dotarray[55][119], dotarray[56][119], dotarray[57][119], dotarray[58][119], dotarray[59][119], dotarray[60][119], dotarray[61][119], dotarray[62][119], dotarray[63][119], dotarray[64][119], dotarray[65][119], dotarray[66][119], dotarray[67][119], dotarray[68][119], dotarray[69][119], dotarray[70][119], dotarray[71][119], dotarray[72][119], dotarray[73][119], dotarray[74][119], dotarray[75][119], dotarray[76][119], dotarray[77][119], dotarray[78][119], dotarray[79][119], dotarray[80][119], dotarray[81][119], dotarray[82][119], dotarray[83][119], dotarray[84][119], dotarray[85][119], dotarray[86][119], dotarray[87][119], dotarray[88][119], dotarray[89][119], dotarray[90][119], dotarray[91][119], dotarray[92][119], dotarray[93][119], dotarray[94][119], dotarray[95][119], dotarray[96][119], dotarray[97][119], dotarray[98][119], dotarray[99][119], dotarray[100][119], dotarray[101][119], dotarray[102][119], dotarray[103][119], dotarray[104][119], dotarray[105][119], dotarray[106][119], dotarray[107][119], dotarray[108][119], dotarray[109][119], dotarray[110][119], dotarray[111][119], dotarray[112][119], dotarray[113][119], dotarray[114][119], dotarray[115][119], dotarray[116][119], dotarray[117][119], dotarray[118][119], dotarray[119][119], dotarray[120][119], dotarray[121][119], dotarray[122][119], dotarray[123][119], dotarray[124][119], dotarray[125][119], dotarray[126][119], dotarray[127][119]};
assign dot_col_120 = {dotarray[0][120], dotarray[1][120], dotarray[2][120], dotarray[3][120], dotarray[4][120], dotarray[5][120], dotarray[6][120], dotarray[7][120], dotarray[8][120], dotarray[9][120], dotarray[10][120], dotarray[11][120], dotarray[12][120], dotarray[13][120], dotarray[14][120], dotarray[15][120], dotarray[16][120], dotarray[17][120], dotarray[18][120], dotarray[19][120], dotarray[20][120], dotarray[21][120], dotarray[22][120], dotarray[23][120], dotarray[24][120], dotarray[25][120], dotarray[26][120], dotarray[27][120], dotarray[28][120], dotarray[29][120], dotarray[30][120], dotarray[31][120], dotarray[32][120], dotarray[33][120], dotarray[34][120], dotarray[35][120], dotarray[36][120], dotarray[37][120], dotarray[38][120], dotarray[39][120], dotarray[40][120], dotarray[41][120], dotarray[42][120], dotarray[43][120], dotarray[44][120], dotarray[45][120], dotarray[46][120], dotarray[47][120], dotarray[48][120], dotarray[49][120], dotarray[50][120], dotarray[51][120], dotarray[52][120], dotarray[53][120], dotarray[54][120], dotarray[55][120], dotarray[56][120], dotarray[57][120], dotarray[58][120], dotarray[59][120], dotarray[60][120], dotarray[61][120], dotarray[62][120], dotarray[63][120], dotarray[64][120], dotarray[65][120], dotarray[66][120], dotarray[67][120], dotarray[68][120], dotarray[69][120], dotarray[70][120], dotarray[71][120], dotarray[72][120], dotarray[73][120], dotarray[74][120], dotarray[75][120], dotarray[76][120], dotarray[77][120], dotarray[78][120], dotarray[79][120], dotarray[80][120], dotarray[81][120], dotarray[82][120], dotarray[83][120], dotarray[84][120], dotarray[85][120], dotarray[86][120], dotarray[87][120], dotarray[88][120], dotarray[89][120], dotarray[90][120], dotarray[91][120], dotarray[92][120], dotarray[93][120], dotarray[94][120], dotarray[95][120], dotarray[96][120], dotarray[97][120], dotarray[98][120], dotarray[99][120], dotarray[100][120], dotarray[101][120], dotarray[102][120], dotarray[103][120], dotarray[104][120], dotarray[105][120], dotarray[106][120], dotarray[107][120], dotarray[108][120], dotarray[109][120], dotarray[110][120], dotarray[111][120], dotarray[112][120], dotarray[113][120], dotarray[114][120], dotarray[115][120], dotarray[116][120], dotarray[117][120], dotarray[118][120], dotarray[119][120], dotarray[120][120], dotarray[121][120], dotarray[122][120], dotarray[123][120], dotarray[124][120], dotarray[125][120], dotarray[126][120], dotarray[127][120]};
assign dot_col_121 = {dotarray[0][121], dotarray[1][121], dotarray[2][121], dotarray[3][121], dotarray[4][121], dotarray[5][121], dotarray[6][121], dotarray[7][121], dotarray[8][121], dotarray[9][121], dotarray[10][121], dotarray[11][121], dotarray[12][121], dotarray[13][121], dotarray[14][121], dotarray[15][121], dotarray[16][121], dotarray[17][121], dotarray[18][121], dotarray[19][121], dotarray[20][121], dotarray[21][121], dotarray[22][121], dotarray[23][121], dotarray[24][121], dotarray[25][121], dotarray[26][121], dotarray[27][121], dotarray[28][121], dotarray[29][121], dotarray[30][121], dotarray[31][121], dotarray[32][121], dotarray[33][121], dotarray[34][121], dotarray[35][121], dotarray[36][121], dotarray[37][121], dotarray[38][121], dotarray[39][121], dotarray[40][121], dotarray[41][121], dotarray[42][121], dotarray[43][121], dotarray[44][121], dotarray[45][121], dotarray[46][121], dotarray[47][121], dotarray[48][121], dotarray[49][121], dotarray[50][121], dotarray[51][121], dotarray[52][121], dotarray[53][121], dotarray[54][121], dotarray[55][121], dotarray[56][121], dotarray[57][121], dotarray[58][121], dotarray[59][121], dotarray[60][121], dotarray[61][121], dotarray[62][121], dotarray[63][121], dotarray[64][121], dotarray[65][121], dotarray[66][121], dotarray[67][121], dotarray[68][121], dotarray[69][121], dotarray[70][121], dotarray[71][121], dotarray[72][121], dotarray[73][121], dotarray[74][121], dotarray[75][121], dotarray[76][121], dotarray[77][121], dotarray[78][121], dotarray[79][121], dotarray[80][121], dotarray[81][121], dotarray[82][121], dotarray[83][121], dotarray[84][121], dotarray[85][121], dotarray[86][121], dotarray[87][121], dotarray[88][121], dotarray[89][121], dotarray[90][121], dotarray[91][121], dotarray[92][121], dotarray[93][121], dotarray[94][121], dotarray[95][121], dotarray[96][121], dotarray[97][121], dotarray[98][121], dotarray[99][121], dotarray[100][121], dotarray[101][121], dotarray[102][121], dotarray[103][121], dotarray[104][121], dotarray[105][121], dotarray[106][121], dotarray[107][121], dotarray[108][121], dotarray[109][121], dotarray[110][121], dotarray[111][121], dotarray[112][121], dotarray[113][121], dotarray[114][121], dotarray[115][121], dotarray[116][121], dotarray[117][121], dotarray[118][121], dotarray[119][121], dotarray[120][121], dotarray[121][121], dotarray[122][121], dotarray[123][121], dotarray[124][121], dotarray[125][121], dotarray[126][121], dotarray[127][121]};
assign dot_col_122 = {dotarray[0][122], dotarray[1][122], dotarray[2][122], dotarray[3][122], dotarray[4][122], dotarray[5][122], dotarray[6][122], dotarray[7][122], dotarray[8][122], dotarray[9][122], dotarray[10][122], dotarray[11][122], dotarray[12][122], dotarray[13][122], dotarray[14][122], dotarray[15][122], dotarray[16][122], dotarray[17][122], dotarray[18][122], dotarray[19][122], dotarray[20][122], dotarray[21][122], dotarray[22][122], dotarray[23][122], dotarray[24][122], dotarray[25][122], dotarray[26][122], dotarray[27][122], dotarray[28][122], dotarray[29][122], dotarray[30][122], dotarray[31][122], dotarray[32][122], dotarray[33][122], dotarray[34][122], dotarray[35][122], dotarray[36][122], dotarray[37][122], dotarray[38][122], dotarray[39][122], dotarray[40][122], dotarray[41][122], dotarray[42][122], dotarray[43][122], dotarray[44][122], dotarray[45][122], dotarray[46][122], dotarray[47][122], dotarray[48][122], dotarray[49][122], dotarray[50][122], dotarray[51][122], dotarray[52][122], dotarray[53][122], dotarray[54][122], dotarray[55][122], dotarray[56][122], dotarray[57][122], dotarray[58][122], dotarray[59][122], dotarray[60][122], dotarray[61][122], dotarray[62][122], dotarray[63][122], dotarray[64][122], dotarray[65][122], dotarray[66][122], dotarray[67][122], dotarray[68][122], dotarray[69][122], dotarray[70][122], dotarray[71][122], dotarray[72][122], dotarray[73][122], dotarray[74][122], dotarray[75][122], dotarray[76][122], dotarray[77][122], dotarray[78][122], dotarray[79][122], dotarray[80][122], dotarray[81][122], dotarray[82][122], dotarray[83][122], dotarray[84][122], dotarray[85][122], dotarray[86][122], dotarray[87][122], dotarray[88][122], dotarray[89][122], dotarray[90][122], dotarray[91][122], dotarray[92][122], dotarray[93][122], dotarray[94][122], dotarray[95][122], dotarray[96][122], dotarray[97][122], dotarray[98][122], dotarray[99][122], dotarray[100][122], dotarray[101][122], dotarray[102][122], dotarray[103][122], dotarray[104][122], dotarray[105][122], dotarray[106][122], dotarray[107][122], dotarray[108][122], dotarray[109][122], dotarray[110][122], dotarray[111][122], dotarray[112][122], dotarray[113][122], dotarray[114][122], dotarray[115][122], dotarray[116][122], dotarray[117][122], dotarray[118][122], dotarray[119][122], dotarray[120][122], dotarray[121][122], dotarray[122][122], dotarray[123][122], dotarray[124][122], dotarray[125][122], dotarray[126][122], dotarray[127][122]};
assign dot_col_123 = {dotarray[0][123], dotarray[1][123], dotarray[2][123], dotarray[3][123], dotarray[4][123], dotarray[5][123], dotarray[6][123], dotarray[7][123], dotarray[8][123], dotarray[9][123], dotarray[10][123], dotarray[11][123], dotarray[12][123], dotarray[13][123], dotarray[14][123], dotarray[15][123], dotarray[16][123], dotarray[17][123], dotarray[18][123], dotarray[19][123], dotarray[20][123], dotarray[21][123], dotarray[22][123], dotarray[23][123], dotarray[24][123], dotarray[25][123], dotarray[26][123], dotarray[27][123], dotarray[28][123], dotarray[29][123], dotarray[30][123], dotarray[31][123], dotarray[32][123], dotarray[33][123], dotarray[34][123], dotarray[35][123], dotarray[36][123], dotarray[37][123], dotarray[38][123], dotarray[39][123], dotarray[40][123], dotarray[41][123], dotarray[42][123], dotarray[43][123], dotarray[44][123], dotarray[45][123], dotarray[46][123], dotarray[47][123], dotarray[48][123], dotarray[49][123], dotarray[50][123], dotarray[51][123], dotarray[52][123], dotarray[53][123], dotarray[54][123], dotarray[55][123], dotarray[56][123], dotarray[57][123], dotarray[58][123], dotarray[59][123], dotarray[60][123], dotarray[61][123], dotarray[62][123], dotarray[63][123], dotarray[64][123], dotarray[65][123], dotarray[66][123], dotarray[67][123], dotarray[68][123], dotarray[69][123], dotarray[70][123], dotarray[71][123], dotarray[72][123], dotarray[73][123], dotarray[74][123], dotarray[75][123], dotarray[76][123], dotarray[77][123], dotarray[78][123], dotarray[79][123], dotarray[80][123], dotarray[81][123], dotarray[82][123], dotarray[83][123], dotarray[84][123], dotarray[85][123], dotarray[86][123], dotarray[87][123], dotarray[88][123], dotarray[89][123], dotarray[90][123], dotarray[91][123], dotarray[92][123], dotarray[93][123], dotarray[94][123], dotarray[95][123], dotarray[96][123], dotarray[97][123], dotarray[98][123], dotarray[99][123], dotarray[100][123], dotarray[101][123], dotarray[102][123], dotarray[103][123], dotarray[104][123], dotarray[105][123], dotarray[106][123], dotarray[107][123], dotarray[108][123], dotarray[109][123], dotarray[110][123], dotarray[111][123], dotarray[112][123], dotarray[113][123], dotarray[114][123], dotarray[115][123], dotarray[116][123], dotarray[117][123], dotarray[118][123], dotarray[119][123], dotarray[120][123], dotarray[121][123], dotarray[122][123], dotarray[123][123], dotarray[124][123], dotarray[125][123], dotarray[126][123], dotarray[127][123]};
assign dot_col_124 = {dotarray[0][124], dotarray[1][124], dotarray[2][124], dotarray[3][124], dotarray[4][124], dotarray[5][124], dotarray[6][124], dotarray[7][124], dotarray[8][124], dotarray[9][124], dotarray[10][124], dotarray[11][124], dotarray[12][124], dotarray[13][124], dotarray[14][124], dotarray[15][124], dotarray[16][124], dotarray[17][124], dotarray[18][124], dotarray[19][124], dotarray[20][124], dotarray[21][124], dotarray[22][124], dotarray[23][124], dotarray[24][124], dotarray[25][124], dotarray[26][124], dotarray[27][124], dotarray[28][124], dotarray[29][124], dotarray[30][124], dotarray[31][124], dotarray[32][124], dotarray[33][124], dotarray[34][124], dotarray[35][124], dotarray[36][124], dotarray[37][124], dotarray[38][124], dotarray[39][124], dotarray[40][124], dotarray[41][124], dotarray[42][124], dotarray[43][124], dotarray[44][124], dotarray[45][124], dotarray[46][124], dotarray[47][124], dotarray[48][124], dotarray[49][124], dotarray[50][124], dotarray[51][124], dotarray[52][124], dotarray[53][124], dotarray[54][124], dotarray[55][124], dotarray[56][124], dotarray[57][124], dotarray[58][124], dotarray[59][124], dotarray[60][124], dotarray[61][124], dotarray[62][124], dotarray[63][124], dotarray[64][124], dotarray[65][124], dotarray[66][124], dotarray[67][124], dotarray[68][124], dotarray[69][124], dotarray[70][124], dotarray[71][124], dotarray[72][124], dotarray[73][124], dotarray[74][124], dotarray[75][124], dotarray[76][124], dotarray[77][124], dotarray[78][124], dotarray[79][124], dotarray[80][124], dotarray[81][124], dotarray[82][124], dotarray[83][124], dotarray[84][124], dotarray[85][124], dotarray[86][124], dotarray[87][124], dotarray[88][124], dotarray[89][124], dotarray[90][124], dotarray[91][124], dotarray[92][124], dotarray[93][124], dotarray[94][124], dotarray[95][124], dotarray[96][124], dotarray[97][124], dotarray[98][124], dotarray[99][124], dotarray[100][124], dotarray[101][124], dotarray[102][124], dotarray[103][124], dotarray[104][124], dotarray[105][124], dotarray[106][124], dotarray[107][124], dotarray[108][124], dotarray[109][124], dotarray[110][124], dotarray[111][124], dotarray[112][124], dotarray[113][124], dotarray[114][124], dotarray[115][124], dotarray[116][124], dotarray[117][124], dotarray[118][124], dotarray[119][124], dotarray[120][124], dotarray[121][124], dotarray[122][124], dotarray[123][124], dotarray[124][124], dotarray[125][124], dotarray[126][124], dotarray[127][124]};
assign dot_col_125 = {dotarray[0][125], dotarray[1][125], dotarray[2][125], dotarray[3][125], dotarray[4][125], dotarray[5][125], dotarray[6][125], dotarray[7][125], dotarray[8][125], dotarray[9][125], dotarray[10][125], dotarray[11][125], dotarray[12][125], dotarray[13][125], dotarray[14][125], dotarray[15][125], dotarray[16][125], dotarray[17][125], dotarray[18][125], dotarray[19][125], dotarray[20][125], dotarray[21][125], dotarray[22][125], dotarray[23][125], dotarray[24][125], dotarray[25][125], dotarray[26][125], dotarray[27][125], dotarray[28][125], dotarray[29][125], dotarray[30][125], dotarray[31][125], dotarray[32][125], dotarray[33][125], dotarray[34][125], dotarray[35][125], dotarray[36][125], dotarray[37][125], dotarray[38][125], dotarray[39][125], dotarray[40][125], dotarray[41][125], dotarray[42][125], dotarray[43][125], dotarray[44][125], dotarray[45][125], dotarray[46][125], dotarray[47][125], dotarray[48][125], dotarray[49][125], dotarray[50][125], dotarray[51][125], dotarray[52][125], dotarray[53][125], dotarray[54][125], dotarray[55][125], dotarray[56][125], dotarray[57][125], dotarray[58][125], dotarray[59][125], dotarray[60][125], dotarray[61][125], dotarray[62][125], dotarray[63][125], dotarray[64][125], dotarray[65][125], dotarray[66][125], dotarray[67][125], dotarray[68][125], dotarray[69][125], dotarray[70][125], dotarray[71][125], dotarray[72][125], dotarray[73][125], dotarray[74][125], dotarray[75][125], dotarray[76][125], dotarray[77][125], dotarray[78][125], dotarray[79][125], dotarray[80][125], dotarray[81][125], dotarray[82][125], dotarray[83][125], dotarray[84][125], dotarray[85][125], dotarray[86][125], dotarray[87][125], dotarray[88][125], dotarray[89][125], dotarray[90][125], dotarray[91][125], dotarray[92][125], dotarray[93][125], dotarray[94][125], dotarray[95][125], dotarray[96][125], dotarray[97][125], dotarray[98][125], dotarray[99][125], dotarray[100][125], dotarray[101][125], dotarray[102][125], dotarray[103][125], dotarray[104][125], dotarray[105][125], dotarray[106][125], dotarray[107][125], dotarray[108][125], dotarray[109][125], dotarray[110][125], dotarray[111][125], dotarray[112][125], dotarray[113][125], dotarray[114][125], dotarray[115][125], dotarray[116][125], dotarray[117][125], dotarray[118][125], dotarray[119][125], dotarray[120][125], dotarray[121][125], dotarray[122][125], dotarray[123][125], dotarray[124][125], dotarray[125][125], dotarray[126][125], dotarray[127][125]};
assign dot_col_126 = {dotarray[0][126], dotarray[1][126], dotarray[2][126], dotarray[3][126], dotarray[4][126], dotarray[5][126], dotarray[6][126], dotarray[7][126], dotarray[8][126], dotarray[9][126], dotarray[10][126], dotarray[11][126], dotarray[12][126], dotarray[13][126], dotarray[14][126], dotarray[15][126], dotarray[16][126], dotarray[17][126], dotarray[18][126], dotarray[19][126], dotarray[20][126], dotarray[21][126], dotarray[22][126], dotarray[23][126], dotarray[24][126], dotarray[25][126], dotarray[26][126], dotarray[27][126], dotarray[28][126], dotarray[29][126], dotarray[30][126], dotarray[31][126], dotarray[32][126], dotarray[33][126], dotarray[34][126], dotarray[35][126], dotarray[36][126], dotarray[37][126], dotarray[38][126], dotarray[39][126], dotarray[40][126], dotarray[41][126], dotarray[42][126], dotarray[43][126], dotarray[44][126], dotarray[45][126], dotarray[46][126], dotarray[47][126], dotarray[48][126], dotarray[49][126], dotarray[50][126], dotarray[51][126], dotarray[52][126], dotarray[53][126], dotarray[54][126], dotarray[55][126], dotarray[56][126], dotarray[57][126], dotarray[58][126], dotarray[59][126], dotarray[60][126], dotarray[61][126], dotarray[62][126], dotarray[63][126], dotarray[64][126], dotarray[65][126], dotarray[66][126], dotarray[67][126], dotarray[68][126], dotarray[69][126], dotarray[70][126], dotarray[71][126], dotarray[72][126], dotarray[73][126], dotarray[74][126], dotarray[75][126], dotarray[76][126], dotarray[77][126], dotarray[78][126], dotarray[79][126], dotarray[80][126], dotarray[81][126], dotarray[82][126], dotarray[83][126], dotarray[84][126], dotarray[85][126], dotarray[86][126], dotarray[87][126], dotarray[88][126], dotarray[89][126], dotarray[90][126], dotarray[91][126], dotarray[92][126], dotarray[93][126], dotarray[94][126], dotarray[95][126], dotarray[96][126], dotarray[97][126], dotarray[98][126], dotarray[99][126], dotarray[100][126], dotarray[101][126], dotarray[102][126], dotarray[103][126], dotarray[104][126], dotarray[105][126], dotarray[106][126], dotarray[107][126], dotarray[108][126], dotarray[109][126], dotarray[110][126], dotarray[111][126], dotarray[112][126], dotarray[113][126], dotarray[114][126], dotarray[115][126], dotarray[116][126], dotarray[117][126], dotarray[118][126], dotarray[119][126], dotarray[120][126], dotarray[121][126], dotarray[122][126], dotarray[123][126], dotarray[124][126], dotarray[125][126], dotarray[126][126], dotarray[127][126]};
assign dot_col_127 = {dotarray[0][127], dotarray[1][127], dotarray[2][127], dotarray[3][127], dotarray[4][127], dotarray[5][127], dotarray[6][127], dotarray[7][127], dotarray[8][127], dotarray[9][127], dotarray[10][127], dotarray[11][127], dotarray[12][127], dotarray[13][127], dotarray[14][127], dotarray[15][127], dotarray[16][127], dotarray[17][127], dotarray[18][127], dotarray[19][127], dotarray[20][127], dotarray[21][127], dotarray[22][127], dotarray[23][127], dotarray[24][127], dotarray[25][127], dotarray[26][127], dotarray[27][127], dotarray[28][127], dotarray[29][127], dotarray[30][127], dotarray[31][127], dotarray[32][127], dotarray[33][127], dotarray[34][127], dotarray[35][127], dotarray[36][127], dotarray[37][127], dotarray[38][127], dotarray[39][127], dotarray[40][127], dotarray[41][127], dotarray[42][127], dotarray[43][127], dotarray[44][127], dotarray[45][127], dotarray[46][127], dotarray[47][127], dotarray[48][127], dotarray[49][127], dotarray[50][127], dotarray[51][127], dotarray[52][127], dotarray[53][127], dotarray[54][127], dotarray[55][127], dotarray[56][127], dotarray[57][127], dotarray[58][127], dotarray[59][127], dotarray[60][127], dotarray[61][127], dotarray[62][127], dotarray[63][127], dotarray[64][127], dotarray[65][127], dotarray[66][127], dotarray[67][127], dotarray[68][127], dotarray[69][127], dotarray[70][127], dotarray[71][127], dotarray[72][127], dotarray[73][127], dotarray[74][127], dotarray[75][127], dotarray[76][127], dotarray[77][127], dotarray[78][127], dotarray[79][127], dotarray[80][127], dotarray[81][127], dotarray[82][127], dotarray[83][127], dotarray[84][127], dotarray[85][127], dotarray[86][127], dotarray[87][127], dotarray[88][127], dotarray[89][127], dotarray[90][127], dotarray[91][127], dotarray[92][127], dotarray[93][127], dotarray[94][127], dotarray[95][127], dotarray[96][127], dotarray[97][127], dotarray[98][127], dotarray[99][127], dotarray[100][127], dotarray[101][127], dotarray[102][127], dotarray[103][127], dotarray[104][127], dotarray[105][127], dotarray[106][127], dotarray[107][127], dotarray[108][127], dotarray[109][127], dotarray[110][127], dotarray[111][127], dotarray[112][127], dotarray[113][127], dotarray[114][127], dotarray[115][127], dotarray[116][127], dotarray[117][127], dotarray[118][127], dotarray[119][127], dotarray[120][127], dotarray[121][127], dotarray[122][127], dotarray[123][127], dotarray[124][127], dotarray[125][127], dotarray[126][127], dotarray[127][127]};
assign dot_col_128 = {dotarray[0][128], dotarray[1][128], dotarray[2][128], dotarray[3][128], dotarray[4][128], dotarray[5][128], dotarray[6][128], dotarray[7][128], dotarray[8][128], dotarray[9][128], dotarray[10][128], dotarray[11][128], dotarray[12][128], dotarray[13][128], dotarray[14][128], dotarray[15][128], dotarray[16][128], dotarray[17][128], dotarray[18][128], dotarray[19][128], dotarray[20][128], dotarray[21][128], dotarray[22][128], dotarray[23][128], dotarray[24][128], dotarray[25][128], dotarray[26][128], dotarray[27][128], dotarray[28][128], dotarray[29][128], dotarray[30][128], dotarray[31][128], dotarray[32][128], dotarray[33][128], dotarray[34][128], dotarray[35][128], dotarray[36][128], dotarray[37][128], dotarray[38][128], dotarray[39][128], dotarray[40][128], dotarray[41][128], dotarray[42][128], dotarray[43][128], dotarray[44][128], dotarray[45][128], dotarray[46][128], dotarray[47][128], dotarray[48][128], dotarray[49][128], dotarray[50][128], dotarray[51][128], dotarray[52][128], dotarray[53][128], dotarray[54][128], dotarray[55][128], dotarray[56][128], dotarray[57][128], dotarray[58][128], dotarray[59][128], dotarray[60][128], dotarray[61][128], dotarray[62][128], dotarray[63][128], dotarray[64][128], dotarray[65][128], dotarray[66][128], dotarray[67][128], dotarray[68][128], dotarray[69][128], dotarray[70][128], dotarray[71][128], dotarray[72][128], dotarray[73][128], dotarray[74][128], dotarray[75][128], dotarray[76][128], dotarray[77][128], dotarray[78][128], dotarray[79][128], dotarray[80][128], dotarray[81][128], dotarray[82][128], dotarray[83][128], dotarray[84][128], dotarray[85][128], dotarray[86][128], dotarray[87][128], dotarray[88][128], dotarray[89][128], dotarray[90][128], dotarray[91][128], dotarray[92][128], dotarray[93][128], dotarray[94][128], dotarray[95][128], dotarray[96][128], dotarray[97][128], dotarray[98][128], dotarray[99][128], dotarray[100][128], dotarray[101][128], dotarray[102][128], dotarray[103][128], dotarray[104][128], dotarray[105][128], dotarray[106][128], dotarray[107][128], dotarray[108][128], dotarray[109][128], dotarray[110][128], dotarray[111][128], dotarray[112][128], dotarray[113][128], dotarray[114][128], dotarray[115][128], dotarray[116][128], dotarray[117][128], dotarray[118][128], dotarray[119][128], dotarray[120][128], dotarray[121][128], dotarray[122][128], dotarray[123][128], dotarray[124][128], dotarray[125][128], dotarray[126][128], dotarray[127][128]};
assign dot_col_129 = {dotarray[0][129], dotarray[1][129], dotarray[2][129], dotarray[3][129], dotarray[4][129], dotarray[5][129], dotarray[6][129], dotarray[7][129], dotarray[8][129], dotarray[9][129], dotarray[10][129], dotarray[11][129], dotarray[12][129], dotarray[13][129], dotarray[14][129], dotarray[15][129], dotarray[16][129], dotarray[17][129], dotarray[18][129], dotarray[19][129], dotarray[20][129], dotarray[21][129], dotarray[22][129], dotarray[23][129], dotarray[24][129], dotarray[25][129], dotarray[26][129], dotarray[27][129], dotarray[28][129], dotarray[29][129], dotarray[30][129], dotarray[31][129], dotarray[32][129], dotarray[33][129], dotarray[34][129], dotarray[35][129], dotarray[36][129], dotarray[37][129], dotarray[38][129], dotarray[39][129], dotarray[40][129], dotarray[41][129], dotarray[42][129], dotarray[43][129], dotarray[44][129], dotarray[45][129], dotarray[46][129], dotarray[47][129], dotarray[48][129], dotarray[49][129], dotarray[50][129], dotarray[51][129], dotarray[52][129], dotarray[53][129], dotarray[54][129], dotarray[55][129], dotarray[56][129], dotarray[57][129], dotarray[58][129], dotarray[59][129], dotarray[60][129], dotarray[61][129], dotarray[62][129], dotarray[63][129], dotarray[64][129], dotarray[65][129], dotarray[66][129], dotarray[67][129], dotarray[68][129], dotarray[69][129], dotarray[70][129], dotarray[71][129], dotarray[72][129], dotarray[73][129], dotarray[74][129], dotarray[75][129], dotarray[76][129], dotarray[77][129], dotarray[78][129], dotarray[79][129], dotarray[80][129], dotarray[81][129], dotarray[82][129], dotarray[83][129], dotarray[84][129], dotarray[85][129], dotarray[86][129], dotarray[87][129], dotarray[88][129], dotarray[89][129], dotarray[90][129], dotarray[91][129], dotarray[92][129], dotarray[93][129], dotarray[94][129], dotarray[95][129], dotarray[96][129], dotarray[97][129], dotarray[98][129], dotarray[99][129], dotarray[100][129], dotarray[101][129], dotarray[102][129], dotarray[103][129], dotarray[104][129], dotarray[105][129], dotarray[106][129], dotarray[107][129], dotarray[108][129], dotarray[109][129], dotarray[110][129], dotarray[111][129], dotarray[112][129], dotarray[113][129], dotarray[114][129], dotarray[115][129], dotarray[116][129], dotarray[117][129], dotarray[118][129], dotarray[119][129], dotarray[120][129], dotarray[121][129], dotarray[122][129], dotarray[123][129], dotarray[124][129], dotarray[125][129], dotarray[126][129], dotarray[127][129]};
assign dot_col_130 = {dotarray[0][130], dotarray[1][130], dotarray[2][130], dotarray[3][130], dotarray[4][130], dotarray[5][130], dotarray[6][130], dotarray[7][130], dotarray[8][130], dotarray[9][130], dotarray[10][130], dotarray[11][130], dotarray[12][130], dotarray[13][130], dotarray[14][130], dotarray[15][130], dotarray[16][130], dotarray[17][130], dotarray[18][130], dotarray[19][130], dotarray[20][130], dotarray[21][130], dotarray[22][130], dotarray[23][130], dotarray[24][130], dotarray[25][130], dotarray[26][130], dotarray[27][130], dotarray[28][130], dotarray[29][130], dotarray[30][130], dotarray[31][130], dotarray[32][130], dotarray[33][130], dotarray[34][130], dotarray[35][130], dotarray[36][130], dotarray[37][130], dotarray[38][130], dotarray[39][130], dotarray[40][130], dotarray[41][130], dotarray[42][130], dotarray[43][130], dotarray[44][130], dotarray[45][130], dotarray[46][130], dotarray[47][130], dotarray[48][130], dotarray[49][130], dotarray[50][130], dotarray[51][130], dotarray[52][130], dotarray[53][130], dotarray[54][130], dotarray[55][130], dotarray[56][130], dotarray[57][130], dotarray[58][130], dotarray[59][130], dotarray[60][130], dotarray[61][130], dotarray[62][130], dotarray[63][130], dotarray[64][130], dotarray[65][130], dotarray[66][130], dotarray[67][130], dotarray[68][130], dotarray[69][130], dotarray[70][130], dotarray[71][130], dotarray[72][130], dotarray[73][130], dotarray[74][130], dotarray[75][130], dotarray[76][130], dotarray[77][130], dotarray[78][130], dotarray[79][130], dotarray[80][130], dotarray[81][130], dotarray[82][130], dotarray[83][130], dotarray[84][130], dotarray[85][130], dotarray[86][130], dotarray[87][130], dotarray[88][130], dotarray[89][130], dotarray[90][130], dotarray[91][130], dotarray[92][130], dotarray[93][130], dotarray[94][130], dotarray[95][130], dotarray[96][130], dotarray[97][130], dotarray[98][130], dotarray[99][130], dotarray[100][130], dotarray[101][130], dotarray[102][130], dotarray[103][130], dotarray[104][130], dotarray[105][130], dotarray[106][130], dotarray[107][130], dotarray[108][130], dotarray[109][130], dotarray[110][130], dotarray[111][130], dotarray[112][130], dotarray[113][130], dotarray[114][130], dotarray[115][130], dotarray[116][130], dotarray[117][130], dotarray[118][130], dotarray[119][130], dotarray[120][130], dotarray[121][130], dotarray[122][130], dotarray[123][130], dotarray[124][130], dotarray[125][130], dotarray[126][130], dotarray[127][130]};
assign dot_col_131 = {dotarray[0][131], dotarray[1][131], dotarray[2][131], dotarray[3][131], dotarray[4][131], dotarray[5][131], dotarray[6][131], dotarray[7][131], dotarray[8][131], dotarray[9][131], dotarray[10][131], dotarray[11][131], dotarray[12][131], dotarray[13][131], dotarray[14][131], dotarray[15][131], dotarray[16][131], dotarray[17][131], dotarray[18][131], dotarray[19][131], dotarray[20][131], dotarray[21][131], dotarray[22][131], dotarray[23][131], dotarray[24][131], dotarray[25][131], dotarray[26][131], dotarray[27][131], dotarray[28][131], dotarray[29][131], dotarray[30][131], dotarray[31][131], dotarray[32][131], dotarray[33][131], dotarray[34][131], dotarray[35][131], dotarray[36][131], dotarray[37][131], dotarray[38][131], dotarray[39][131], dotarray[40][131], dotarray[41][131], dotarray[42][131], dotarray[43][131], dotarray[44][131], dotarray[45][131], dotarray[46][131], dotarray[47][131], dotarray[48][131], dotarray[49][131], dotarray[50][131], dotarray[51][131], dotarray[52][131], dotarray[53][131], dotarray[54][131], dotarray[55][131], dotarray[56][131], dotarray[57][131], dotarray[58][131], dotarray[59][131], dotarray[60][131], dotarray[61][131], dotarray[62][131], dotarray[63][131], dotarray[64][131], dotarray[65][131], dotarray[66][131], dotarray[67][131], dotarray[68][131], dotarray[69][131], dotarray[70][131], dotarray[71][131], dotarray[72][131], dotarray[73][131], dotarray[74][131], dotarray[75][131], dotarray[76][131], dotarray[77][131], dotarray[78][131], dotarray[79][131], dotarray[80][131], dotarray[81][131], dotarray[82][131], dotarray[83][131], dotarray[84][131], dotarray[85][131], dotarray[86][131], dotarray[87][131], dotarray[88][131], dotarray[89][131], dotarray[90][131], dotarray[91][131], dotarray[92][131], dotarray[93][131], dotarray[94][131], dotarray[95][131], dotarray[96][131], dotarray[97][131], dotarray[98][131], dotarray[99][131], dotarray[100][131], dotarray[101][131], dotarray[102][131], dotarray[103][131], dotarray[104][131], dotarray[105][131], dotarray[106][131], dotarray[107][131], dotarray[108][131], dotarray[109][131], dotarray[110][131], dotarray[111][131], dotarray[112][131], dotarray[113][131], dotarray[114][131], dotarray[115][131], dotarray[116][131], dotarray[117][131], dotarray[118][131], dotarray[119][131], dotarray[120][131], dotarray[121][131], dotarray[122][131], dotarray[123][131], dotarray[124][131], dotarray[125][131], dotarray[126][131], dotarray[127][131]};
assign dot_col_132 = {dotarray[0][132], dotarray[1][132], dotarray[2][132], dotarray[3][132], dotarray[4][132], dotarray[5][132], dotarray[6][132], dotarray[7][132], dotarray[8][132], dotarray[9][132], dotarray[10][132], dotarray[11][132], dotarray[12][132], dotarray[13][132], dotarray[14][132], dotarray[15][132], dotarray[16][132], dotarray[17][132], dotarray[18][132], dotarray[19][132], dotarray[20][132], dotarray[21][132], dotarray[22][132], dotarray[23][132], dotarray[24][132], dotarray[25][132], dotarray[26][132], dotarray[27][132], dotarray[28][132], dotarray[29][132], dotarray[30][132], dotarray[31][132], dotarray[32][132], dotarray[33][132], dotarray[34][132], dotarray[35][132], dotarray[36][132], dotarray[37][132], dotarray[38][132], dotarray[39][132], dotarray[40][132], dotarray[41][132], dotarray[42][132], dotarray[43][132], dotarray[44][132], dotarray[45][132], dotarray[46][132], dotarray[47][132], dotarray[48][132], dotarray[49][132], dotarray[50][132], dotarray[51][132], dotarray[52][132], dotarray[53][132], dotarray[54][132], dotarray[55][132], dotarray[56][132], dotarray[57][132], dotarray[58][132], dotarray[59][132], dotarray[60][132], dotarray[61][132], dotarray[62][132], dotarray[63][132], dotarray[64][132], dotarray[65][132], dotarray[66][132], dotarray[67][132], dotarray[68][132], dotarray[69][132], dotarray[70][132], dotarray[71][132], dotarray[72][132], dotarray[73][132], dotarray[74][132], dotarray[75][132], dotarray[76][132], dotarray[77][132], dotarray[78][132], dotarray[79][132], dotarray[80][132], dotarray[81][132], dotarray[82][132], dotarray[83][132], dotarray[84][132], dotarray[85][132], dotarray[86][132], dotarray[87][132], dotarray[88][132], dotarray[89][132], dotarray[90][132], dotarray[91][132], dotarray[92][132], dotarray[93][132], dotarray[94][132], dotarray[95][132], dotarray[96][132], dotarray[97][132], dotarray[98][132], dotarray[99][132], dotarray[100][132], dotarray[101][132], dotarray[102][132], dotarray[103][132], dotarray[104][132], dotarray[105][132], dotarray[106][132], dotarray[107][132], dotarray[108][132], dotarray[109][132], dotarray[110][132], dotarray[111][132], dotarray[112][132], dotarray[113][132], dotarray[114][132], dotarray[115][132], dotarray[116][132], dotarray[117][132], dotarray[118][132], dotarray[119][132], dotarray[120][132], dotarray[121][132], dotarray[122][132], dotarray[123][132], dotarray[124][132], dotarray[125][132], dotarray[126][132], dotarray[127][132]};
assign dot_col_133 = {dotarray[0][133], dotarray[1][133], dotarray[2][133], dotarray[3][133], dotarray[4][133], dotarray[5][133], dotarray[6][133], dotarray[7][133], dotarray[8][133], dotarray[9][133], dotarray[10][133], dotarray[11][133], dotarray[12][133], dotarray[13][133], dotarray[14][133], dotarray[15][133], dotarray[16][133], dotarray[17][133], dotarray[18][133], dotarray[19][133], dotarray[20][133], dotarray[21][133], dotarray[22][133], dotarray[23][133], dotarray[24][133], dotarray[25][133], dotarray[26][133], dotarray[27][133], dotarray[28][133], dotarray[29][133], dotarray[30][133], dotarray[31][133], dotarray[32][133], dotarray[33][133], dotarray[34][133], dotarray[35][133], dotarray[36][133], dotarray[37][133], dotarray[38][133], dotarray[39][133], dotarray[40][133], dotarray[41][133], dotarray[42][133], dotarray[43][133], dotarray[44][133], dotarray[45][133], dotarray[46][133], dotarray[47][133], dotarray[48][133], dotarray[49][133], dotarray[50][133], dotarray[51][133], dotarray[52][133], dotarray[53][133], dotarray[54][133], dotarray[55][133], dotarray[56][133], dotarray[57][133], dotarray[58][133], dotarray[59][133], dotarray[60][133], dotarray[61][133], dotarray[62][133], dotarray[63][133], dotarray[64][133], dotarray[65][133], dotarray[66][133], dotarray[67][133], dotarray[68][133], dotarray[69][133], dotarray[70][133], dotarray[71][133], dotarray[72][133], dotarray[73][133], dotarray[74][133], dotarray[75][133], dotarray[76][133], dotarray[77][133], dotarray[78][133], dotarray[79][133], dotarray[80][133], dotarray[81][133], dotarray[82][133], dotarray[83][133], dotarray[84][133], dotarray[85][133], dotarray[86][133], dotarray[87][133], dotarray[88][133], dotarray[89][133], dotarray[90][133], dotarray[91][133], dotarray[92][133], dotarray[93][133], dotarray[94][133], dotarray[95][133], dotarray[96][133], dotarray[97][133], dotarray[98][133], dotarray[99][133], dotarray[100][133], dotarray[101][133], dotarray[102][133], dotarray[103][133], dotarray[104][133], dotarray[105][133], dotarray[106][133], dotarray[107][133], dotarray[108][133], dotarray[109][133], dotarray[110][133], dotarray[111][133], dotarray[112][133], dotarray[113][133], dotarray[114][133], dotarray[115][133], dotarray[116][133], dotarray[117][133], dotarray[118][133], dotarray[119][133], dotarray[120][133], dotarray[121][133], dotarray[122][133], dotarray[123][133], dotarray[124][133], dotarray[125][133], dotarray[126][133], dotarray[127][133]};
assign dot_col_134 = {dotarray[0][134], dotarray[1][134], dotarray[2][134], dotarray[3][134], dotarray[4][134], dotarray[5][134], dotarray[6][134], dotarray[7][134], dotarray[8][134], dotarray[9][134], dotarray[10][134], dotarray[11][134], dotarray[12][134], dotarray[13][134], dotarray[14][134], dotarray[15][134], dotarray[16][134], dotarray[17][134], dotarray[18][134], dotarray[19][134], dotarray[20][134], dotarray[21][134], dotarray[22][134], dotarray[23][134], dotarray[24][134], dotarray[25][134], dotarray[26][134], dotarray[27][134], dotarray[28][134], dotarray[29][134], dotarray[30][134], dotarray[31][134], dotarray[32][134], dotarray[33][134], dotarray[34][134], dotarray[35][134], dotarray[36][134], dotarray[37][134], dotarray[38][134], dotarray[39][134], dotarray[40][134], dotarray[41][134], dotarray[42][134], dotarray[43][134], dotarray[44][134], dotarray[45][134], dotarray[46][134], dotarray[47][134], dotarray[48][134], dotarray[49][134], dotarray[50][134], dotarray[51][134], dotarray[52][134], dotarray[53][134], dotarray[54][134], dotarray[55][134], dotarray[56][134], dotarray[57][134], dotarray[58][134], dotarray[59][134], dotarray[60][134], dotarray[61][134], dotarray[62][134], dotarray[63][134], dotarray[64][134], dotarray[65][134], dotarray[66][134], dotarray[67][134], dotarray[68][134], dotarray[69][134], dotarray[70][134], dotarray[71][134], dotarray[72][134], dotarray[73][134], dotarray[74][134], dotarray[75][134], dotarray[76][134], dotarray[77][134], dotarray[78][134], dotarray[79][134], dotarray[80][134], dotarray[81][134], dotarray[82][134], dotarray[83][134], dotarray[84][134], dotarray[85][134], dotarray[86][134], dotarray[87][134], dotarray[88][134], dotarray[89][134], dotarray[90][134], dotarray[91][134], dotarray[92][134], dotarray[93][134], dotarray[94][134], dotarray[95][134], dotarray[96][134], dotarray[97][134], dotarray[98][134], dotarray[99][134], dotarray[100][134], dotarray[101][134], dotarray[102][134], dotarray[103][134], dotarray[104][134], dotarray[105][134], dotarray[106][134], dotarray[107][134], dotarray[108][134], dotarray[109][134], dotarray[110][134], dotarray[111][134], dotarray[112][134], dotarray[113][134], dotarray[114][134], dotarray[115][134], dotarray[116][134], dotarray[117][134], dotarray[118][134], dotarray[119][134], dotarray[120][134], dotarray[121][134], dotarray[122][134], dotarray[123][134], dotarray[124][134], dotarray[125][134], dotarray[126][134], dotarray[127][134]};
assign dot_col_135 = {dotarray[0][135], dotarray[1][135], dotarray[2][135], dotarray[3][135], dotarray[4][135], dotarray[5][135], dotarray[6][135], dotarray[7][135], dotarray[8][135], dotarray[9][135], dotarray[10][135], dotarray[11][135], dotarray[12][135], dotarray[13][135], dotarray[14][135], dotarray[15][135], dotarray[16][135], dotarray[17][135], dotarray[18][135], dotarray[19][135], dotarray[20][135], dotarray[21][135], dotarray[22][135], dotarray[23][135], dotarray[24][135], dotarray[25][135], dotarray[26][135], dotarray[27][135], dotarray[28][135], dotarray[29][135], dotarray[30][135], dotarray[31][135], dotarray[32][135], dotarray[33][135], dotarray[34][135], dotarray[35][135], dotarray[36][135], dotarray[37][135], dotarray[38][135], dotarray[39][135], dotarray[40][135], dotarray[41][135], dotarray[42][135], dotarray[43][135], dotarray[44][135], dotarray[45][135], dotarray[46][135], dotarray[47][135], dotarray[48][135], dotarray[49][135], dotarray[50][135], dotarray[51][135], dotarray[52][135], dotarray[53][135], dotarray[54][135], dotarray[55][135], dotarray[56][135], dotarray[57][135], dotarray[58][135], dotarray[59][135], dotarray[60][135], dotarray[61][135], dotarray[62][135], dotarray[63][135], dotarray[64][135], dotarray[65][135], dotarray[66][135], dotarray[67][135], dotarray[68][135], dotarray[69][135], dotarray[70][135], dotarray[71][135], dotarray[72][135], dotarray[73][135], dotarray[74][135], dotarray[75][135], dotarray[76][135], dotarray[77][135], dotarray[78][135], dotarray[79][135], dotarray[80][135], dotarray[81][135], dotarray[82][135], dotarray[83][135], dotarray[84][135], dotarray[85][135], dotarray[86][135], dotarray[87][135], dotarray[88][135], dotarray[89][135], dotarray[90][135], dotarray[91][135], dotarray[92][135], dotarray[93][135], dotarray[94][135], dotarray[95][135], dotarray[96][135], dotarray[97][135], dotarray[98][135], dotarray[99][135], dotarray[100][135], dotarray[101][135], dotarray[102][135], dotarray[103][135], dotarray[104][135], dotarray[105][135], dotarray[106][135], dotarray[107][135], dotarray[108][135], dotarray[109][135], dotarray[110][135], dotarray[111][135], dotarray[112][135], dotarray[113][135], dotarray[114][135], dotarray[115][135], dotarray[116][135], dotarray[117][135], dotarray[118][135], dotarray[119][135], dotarray[120][135], dotarray[121][135], dotarray[122][135], dotarray[123][135], dotarray[124][135], dotarray[125][135], dotarray[126][135], dotarray[127][135]};
assign dot_col_136 = {dotarray[0][136], dotarray[1][136], dotarray[2][136], dotarray[3][136], dotarray[4][136], dotarray[5][136], dotarray[6][136], dotarray[7][136], dotarray[8][136], dotarray[9][136], dotarray[10][136], dotarray[11][136], dotarray[12][136], dotarray[13][136], dotarray[14][136], dotarray[15][136], dotarray[16][136], dotarray[17][136], dotarray[18][136], dotarray[19][136], dotarray[20][136], dotarray[21][136], dotarray[22][136], dotarray[23][136], dotarray[24][136], dotarray[25][136], dotarray[26][136], dotarray[27][136], dotarray[28][136], dotarray[29][136], dotarray[30][136], dotarray[31][136], dotarray[32][136], dotarray[33][136], dotarray[34][136], dotarray[35][136], dotarray[36][136], dotarray[37][136], dotarray[38][136], dotarray[39][136], dotarray[40][136], dotarray[41][136], dotarray[42][136], dotarray[43][136], dotarray[44][136], dotarray[45][136], dotarray[46][136], dotarray[47][136], dotarray[48][136], dotarray[49][136], dotarray[50][136], dotarray[51][136], dotarray[52][136], dotarray[53][136], dotarray[54][136], dotarray[55][136], dotarray[56][136], dotarray[57][136], dotarray[58][136], dotarray[59][136], dotarray[60][136], dotarray[61][136], dotarray[62][136], dotarray[63][136], dotarray[64][136], dotarray[65][136], dotarray[66][136], dotarray[67][136], dotarray[68][136], dotarray[69][136], dotarray[70][136], dotarray[71][136], dotarray[72][136], dotarray[73][136], dotarray[74][136], dotarray[75][136], dotarray[76][136], dotarray[77][136], dotarray[78][136], dotarray[79][136], dotarray[80][136], dotarray[81][136], dotarray[82][136], dotarray[83][136], dotarray[84][136], dotarray[85][136], dotarray[86][136], dotarray[87][136], dotarray[88][136], dotarray[89][136], dotarray[90][136], dotarray[91][136], dotarray[92][136], dotarray[93][136], dotarray[94][136], dotarray[95][136], dotarray[96][136], dotarray[97][136], dotarray[98][136], dotarray[99][136], dotarray[100][136], dotarray[101][136], dotarray[102][136], dotarray[103][136], dotarray[104][136], dotarray[105][136], dotarray[106][136], dotarray[107][136], dotarray[108][136], dotarray[109][136], dotarray[110][136], dotarray[111][136], dotarray[112][136], dotarray[113][136], dotarray[114][136], dotarray[115][136], dotarray[116][136], dotarray[117][136], dotarray[118][136], dotarray[119][136], dotarray[120][136], dotarray[121][136], dotarray[122][136], dotarray[123][136], dotarray[124][136], dotarray[125][136], dotarray[126][136], dotarray[127][136]};
assign dot_col_137 = {dotarray[0][137], dotarray[1][137], dotarray[2][137], dotarray[3][137], dotarray[4][137], dotarray[5][137], dotarray[6][137], dotarray[7][137], dotarray[8][137], dotarray[9][137], dotarray[10][137], dotarray[11][137], dotarray[12][137], dotarray[13][137], dotarray[14][137], dotarray[15][137], dotarray[16][137], dotarray[17][137], dotarray[18][137], dotarray[19][137], dotarray[20][137], dotarray[21][137], dotarray[22][137], dotarray[23][137], dotarray[24][137], dotarray[25][137], dotarray[26][137], dotarray[27][137], dotarray[28][137], dotarray[29][137], dotarray[30][137], dotarray[31][137], dotarray[32][137], dotarray[33][137], dotarray[34][137], dotarray[35][137], dotarray[36][137], dotarray[37][137], dotarray[38][137], dotarray[39][137], dotarray[40][137], dotarray[41][137], dotarray[42][137], dotarray[43][137], dotarray[44][137], dotarray[45][137], dotarray[46][137], dotarray[47][137], dotarray[48][137], dotarray[49][137], dotarray[50][137], dotarray[51][137], dotarray[52][137], dotarray[53][137], dotarray[54][137], dotarray[55][137], dotarray[56][137], dotarray[57][137], dotarray[58][137], dotarray[59][137], dotarray[60][137], dotarray[61][137], dotarray[62][137], dotarray[63][137], dotarray[64][137], dotarray[65][137], dotarray[66][137], dotarray[67][137], dotarray[68][137], dotarray[69][137], dotarray[70][137], dotarray[71][137], dotarray[72][137], dotarray[73][137], dotarray[74][137], dotarray[75][137], dotarray[76][137], dotarray[77][137], dotarray[78][137], dotarray[79][137], dotarray[80][137], dotarray[81][137], dotarray[82][137], dotarray[83][137], dotarray[84][137], dotarray[85][137], dotarray[86][137], dotarray[87][137], dotarray[88][137], dotarray[89][137], dotarray[90][137], dotarray[91][137], dotarray[92][137], dotarray[93][137], dotarray[94][137], dotarray[95][137], dotarray[96][137], dotarray[97][137], dotarray[98][137], dotarray[99][137], dotarray[100][137], dotarray[101][137], dotarray[102][137], dotarray[103][137], dotarray[104][137], dotarray[105][137], dotarray[106][137], dotarray[107][137], dotarray[108][137], dotarray[109][137], dotarray[110][137], dotarray[111][137], dotarray[112][137], dotarray[113][137], dotarray[114][137], dotarray[115][137], dotarray[116][137], dotarray[117][137], dotarray[118][137], dotarray[119][137], dotarray[120][137], dotarray[121][137], dotarray[122][137], dotarray[123][137], dotarray[124][137], dotarray[125][137], dotarray[126][137], dotarray[127][137]};
assign dot_col_138 = {dotarray[0][138], dotarray[1][138], dotarray[2][138], dotarray[3][138], dotarray[4][138], dotarray[5][138], dotarray[6][138], dotarray[7][138], dotarray[8][138], dotarray[9][138], dotarray[10][138], dotarray[11][138], dotarray[12][138], dotarray[13][138], dotarray[14][138], dotarray[15][138], dotarray[16][138], dotarray[17][138], dotarray[18][138], dotarray[19][138], dotarray[20][138], dotarray[21][138], dotarray[22][138], dotarray[23][138], dotarray[24][138], dotarray[25][138], dotarray[26][138], dotarray[27][138], dotarray[28][138], dotarray[29][138], dotarray[30][138], dotarray[31][138], dotarray[32][138], dotarray[33][138], dotarray[34][138], dotarray[35][138], dotarray[36][138], dotarray[37][138], dotarray[38][138], dotarray[39][138], dotarray[40][138], dotarray[41][138], dotarray[42][138], dotarray[43][138], dotarray[44][138], dotarray[45][138], dotarray[46][138], dotarray[47][138], dotarray[48][138], dotarray[49][138], dotarray[50][138], dotarray[51][138], dotarray[52][138], dotarray[53][138], dotarray[54][138], dotarray[55][138], dotarray[56][138], dotarray[57][138], dotarray[58][138], dotarray[59][138], dotarray[60][138], dotarray[61][138], dotarray[62][138], dotarray[63][138], dotarray[64][138], dotarray[65][138], dotarray[66][138], dotarray[67][138], dotarray[68][138], dotarray[69][138], dotarray[70][138], dotarray[71][138], dotarray[72][138], dotarray[73][138], dotarray[74][138], dotarray[75][138], dotarray[76][138], dotarray[77][138], dotarray[78][138], dotarray[79][138], dotarray[80][138], dotarray[81][138], dotarray[82][138], dotarray[83][138], dotarray[84][138], dotarray[85][138], dotarray[86][138], dotarray[87][138], dotarray[88][138], dotarray[89][138], dotarray[90][138], dotarray[91][138], dotarray[92][138], dotarray[93][138], dotarray[94][138], dotarray[95][138], dotarray[96][138], dotarray[97][138], dotarray[98][138], dotarray[99][138], dotarray[100][138], dotarray[101][138], dotarray[102][138], dotarray[103][138], dotarray[104][138], dotarray[105][138], dotarray[106][138], dotarray[107][138], dotarray[108][138], dotarray[109][138], dotarray[110][138], dotarray[111][138], dotarray[112][138], dotarray[113][138], dotarray[114][138], dotarray[115][138], dotarray[116][138], dotarray[117][138], dotarray[118][138], dotarray[119][138], dotarray[120][138], dotarray[121][138], dotarray[122][138], dotarray[123][138], dotarray[124][138], dotarray[125][138], dotarray[126][138], dotarray[127][138]};
assign dot_col_139 = {dotarray[0][139], dotarray[1][139], dotarray[2][139], dotarray[3][139], dotarray[4][139], dotarray[5][139], dotarray[6][139], dotarray[7][139], dotarray[8][139], dotarray[9][139], dotarray[10][139], dotarray[11][139], dotarray[12][139], dotarray[13][139], dotarray[14][139], dotarray[15][139], dotarray[16][139], dotarray[17][139], dotarray[18][139], dotarray[19][139], dotarray[20][139], dotarray[21][139], dotarray[22][139], dotarray[23][139], dotarray[24][139], dotarray[25][139], dotarray[26][139], dotarray[27][139], dotarray[28][139], dotarray[29][139], dotarray[30][139], dotarray[31][139], dotarray[32][139], dotarray[33][139], dotarray[34][139], dotarray[35][139], dotarray[36][139], dotarray[37][139], dotarray[38][139], dotarray[39][139], dotarray[40][139], dotarray[41][139], dotarray[42][139], dotarray[43][139], dotarray[44][139], dotarray[45][139], dotarray[46][139], dotarray[47][139], dotarray[48][139], dotarray[49][139], dotarray[50][139], dotarray[51][139], dotarray[52][139], dotarray[53][139], dotarray[54][139], dotarray[55][139], dotarray[56][139], dotarray[57][139], dotarray[58][139], dotarray[59][139], dotarray[60][139], dotarray[61][139], dotarray[62][139], dotarray[63][139], dotarray[64][139], dotarray[65][139], dotarray[66][139], dotarray[67][139], dotarray[68][139], dotarray[69][139], dotarray[70][139], dotarray[71][139], dotarray[72][139], dotarray[73][139], dotarray[74][139], dotarray[75][139], dotarray[76][139], dotarray[77][139], dotarray[78][139], dotarray[79][139], dotarray[80][139], dotarray[81][139], dotarray[82][139], dotarray[83][139], dotarray[84][139], dotarray[85][139], dotarray[86][139], dotarray[87][139], dotarray[88][139], dotarray[89][139], dotarray[90][139], dotarray[91][139], dotarray[92][139], dotarray[93][139], dotarray[94][139], dotarray[95][139], dotarray[96][139], dotarray[97][139], dotarray[98][139], dotarray[99][139], dotarray[100][139], dotarray[101][139], dotarray[102][139], dotarray[103][139], dotarray[104][139], dotarray[105][139], dotarray[106][139], dotarray[107][139], dotarray[108][139], dotarray[109][139], dotarray[110][139], dotarray[111][139], dotarray[112][139], dotarray[113][139], dotarray[114][139], dotarray[115][139], dotarray[116][139], dotarray[117][139], dotarray[118][139], dotarray[119][139], dotarray[120][139], dotarray[121][139], dotarray[122][139], dotarray[123][139], dotarray[124][139], dotarray[125][139], dotarray[126][139], dotarray[127][139]};
assign dot_col_140 = {dotarray[0][140], dotarray[1][140], dotarray[2][140], dotarray[3][140], dotarray[4][140], dotarray[5][140], dotarray[6][140], dotarray[7][140], dotarray[8][140], dotarray[9][140], dotarray[10][140], dotarray[11][140], dotarray[12][140], dotarray[13][140], dotarray[14][140], dotarray[15][140], dotarray[16][140], dotarray[17][140], dotarray[18][140], dotarray[19][140], dotarray[20][140], dotarray[21][140], dotarray[22][140], dotarray[23][140], dotarray[24][140], dotarray[25][140], dotarray[26][140], dotarray[27][140], dotarray[28][140], dotarray[29][140], dotarray[30][140], dotarray[31][140], dotarray[32][140], dotarray[33][140], dotarray[34][140], dotarray[35][140], dotarray[36][140], dotarray[37][140], dotarray[38][140], dotarray[39][140], dotarray[40][140], dotarray[41][140], dotarray[42][140], dotarray[43][140], dotarray[44][140], dotarray[45][140], dotarray[46][140], dotarray[47][140], dotarray[48][140], dotarray[49][140], dotarray[50][140], dotarray[51][140], dotarray[52][140], dotarray[53][140], dotarray[54][140], dotarray[55][140], dotarray[56][140], dotarray[57][140], dotarray[58][140], dotarray[59][140], dotarray[60][140], dotarray[61][140], dotarray[62][140], dotarray[63][140], dotarray[64][140], dotarray[65][140], dotarray[66][140], dotarray[67][140], dotarray[68][140], dotarray[69][140], dotarray[70][140], dotarray[71][140], dotarray[72][140], dotarray[73][140], dotarray[74][140], dotarray[75][140], dotarray[76][140], dotarray[77][140], dotarray[78][140], dotarray[79][140], dotarray[80][140], dotarray[81][140], dotarray[82][140], dotarray[83][140], dotarray[84][140], dotarray[85][140], dotarray[86][140], dotarray[87][140], dotarray[88][140], dotarray[89][140], dotarray[90][140], dotarray[91][140], dotarray[92][140], dotarray[93][140], dotarray[94][140], dotarray[95][140], dotarray[96][140], dotarray[97][140], dotarray[98][140], dotarray[99][140], dotarray[100][140], dotarray[101][140], dotarray[102][140], dotarray[103][140], dotarray[104][140], dotarray[105][140], dotarray[106][140], dotarray[107][140], dotarray[108][140], dotarray[109][140], dotarray[110][140], dotarray[111][140], dotarray[112][140], dotarray[113][140], dotarray[114][140], dotarray[115][140], dotarray[116][140], dotarray[117][140], dotarray[118][140], dotarray[119][140], dotarray[120][140], dotarray[121][140], dotarray[122][140], dotarray[123][140], dotarray[124][140], dotarray[125][140], dotarray[126][140], dotarray[127][140]};
assign dot_col_141 = {dotarray[0][141], dotarray[1][141], dotarray[2][141], dotarray[3][141], dotarray[4][141], dotarray[5][141], dotarray[6][141], dotarray[7][141], dotarray[8][141], dotarray[9][141], dotarray[10][141], dotarray[11][141], dotarray[12][141], dotarray[13][141], dotarray[14][141], dotarray[15][141], dotarray[16][141], dotarray[17][141], dotarray[18][141], dotarray[19][141], dotarray[20][141], dotarray[21][141], dotarray[22][141], dotarray[23][141], dotarray[24][141], dotarray[25][141], dotarray[26][141], dotarray[27][141], dotarray[28][141], dotarray[29][141], dotarray[30][141], dotarray[31][141], dotarray[32][141], dotarray[33][141], dotarray[34][141], dotarray[35][141], dotarray[36][141], dotarray[37][141], dotarray[38][141], dotarray[39][141], dotarray[40][141], dotarray[41][141], dotarray[42][141], dotarray[43][141], dotarray[44][141], dotarray[45][141], dotarray[46][141], dotarray[47][141], dotarray[48][141], dotarray[49][141], dotarray[50][141], dotarray[51][141], dotarray[52][141], dotarray[53][141], dotarray[54][141], dotarray[55][141], dotarray[56][141], dotarray[57][141], dotarray[58][141], dotarray[59][141], dotarray[60][141], dotarray[61][141], dotarray[62][141], dotarray[63][141], dotarray[64][141], dotarray[65][141], dotarray[66][141], dotarray[67][141], dotarray[68][141], dotarray[69][141], dotarray[70][141], dotarray[71][141], dotarray[72][141], dotarray[73][141], dotarray[74][141], dotarray[75][141], dotarray[76][141], dotarray[77][141], dotarray[78][141], dotarray[79][141], dotarray[80][141], dotarray[81][141], dotarray[82][141], dotarray[83][141], dotarray[84][141], dotarray[85][141], dotarray[86][141], dotarray[87][141], dotarray[88][141], dotarray[89][141], dotarray[90][141], dotarray[91][141], dotarray[92][141], dotarray[93][141], dotarray[94][141], dotarray[95][141], dotarray[96][141], dotarray[97][141], dotarray[98][141], dotarray[99][141], dotarray[100][141], dotarray[101][141], dotarray[102][141], dotarray[103][141], dotarray[104][141], dotarray[105][141], dotarray[106][141], dotarray[107][141], dotarray[108][141], dotarray[109][141], dotarray[110][141], dotarray[111][141], dotarray[112][141], dotarray[113][141], dotarray[114][141], dotarray[115][141], dotarray[116][141], dotarray[117][141], dotarray[118][141], dotarray[119][141], dotarray[120][141], dotarray[121][141], dotarray[122][141], dotarray[123][141], dotarray[124][141], dotarray[125][141], dotarray[126][141], dotarray[127][141]};
assign dot_col_142 = {dotarray[0][142], dotarray[1][142], dotarray[2][142], dotarray[3][142], dotarray[4][142], dotarray[5][142], dotarray[6][142], dotarray[7][142], dotarray[8][142], dotarray[9][142], dotarray[10][142], dotarray[11][142], dotarray[12][142], dotarray[13][142], dotarray[14][142], dotarray[15][142], dotarray[16][142], dotarray[17][142], dotarray[18][142], dotarray[19][142], dotarray[20][142], dotarray[21][142], dotarray[22][142], dotarray[23][142], dotarray[24][142], dotarray[25][142], dotarray[26][142], dotarray[27][142], dotarray[28][142], dotarray[29][142], dotarray[30][142], dotarray[31][142], dotarray[32][142], dotarray[33][142], dotarray[34][142], dotarray[35][142], dotarray[36][142], dotarray[37][142], dotarray[38][142], dotarray[39][142], dotarray[40][142], dotarray[41][142], dotarray[42][142], dotarray[43][142], dotarray[44][142], dotarray[45][142], dotarray[46][142], dotarray[47][142], dotarray[48][142], dotarray[49][142], dotarray[50][142], dotarray[51][142], dotarray[52][142], dotarray[53][142], dotarray[54][142], dotarray[55][142], dotarray[56][142], dotarray[57][142], dotarray[58][142], dotarray[59][142], dotarray[60][142], dotarray[61][142], dotarray[62][142], dotarray[63][142], dotarray[64][142], dotarray[65][142], dotarray[66][142], dotarray[67][142], dotarray[68][142], dotarray[69][142], dotarray[70][142], dotarray[71][142], dotarray[72][142], dotarray[73][142], dotarray[74][142], dotarray[75][142], dotarray[76][142], dotarray[77][142], dotarray[78][142], dotarray[79][142], dotarray[80][142], dotarray[81][142], dotarray[82][142], dotarray[83][142], dotarray[84][142], dotarray[85][142], dotarray[86][142], dotarray[87][142], dotarray[88][142], dotarray[89][142], dotarray[90][142], dotarray[91][142], dotarray[92][142], dotarray[93][142], dotarray[94][142], dotarray[95][142], dotarray[96][142], dotarray[97][142], dotarray[98][142], dotarray[99][142], dotarray[100][142], dotarray[101][142], dotarray[102][142], dotarray[103][142], dotarray[104][142], dotarray[105][142], dotarray[106][142], dotarray[107][142], dotarray[108][142], dotarray[109][142], dotarray[110][142], dotarray[111][142], dotarray[112][142], dotarray[113][142], dotarray[114][142], dotarray[115][142], dotarray[116][142], dotarray[117][142], dotarray[118][142], dotarray[119][142], dotarray[120][142], dotarray[121][142], dotarray[122][142], dotarray[123][142], dotarray[124][142], dotarray[125][142], dotarray[126][142], dotarray[127][142]};
assign dot_col_143 = {dotarray[0][143], dotarray[1][143], dotarray[2][143], dotarray[3][143], dotarray[4][143], dotarray[5][143], dotarray[6][143], dotarray[7][143], dotarray[8][143], dotarray[9][143], dotarray[10][143], dotarray[11][143], dotarray[12][143], dotarray[13][143], dotarray[14][143], dotarray[15][143], dotarray[16][143], dotarray[17][143], dotarray[18][143], dotarray[19][143], dotarray[20][143], dotarray[21][143], dotarray[22][143], dotarray[23][143], dotarray[24][143], dotarray[25][143], dotarray[26][143], dotarray[27][143], dotarray[28][143], dotarray[29][143], dotarray[30][143], dotarray[31][143], dotarray[32][143], dotarray[33][143], dotarray[34][143], dotarray[35][143], dotarray[36][143], dotarray[37][143], dotarray[38][143], dotarray[39][143], dotarray[40][143], dotarray[41][143], dotarray[42][143], dotarray[43][143], dotarray[44][143], dotarray[45][143], dotarray[46][143], dotarray[47][143], dotarray[48][143], dotarray[49][143], dotarray[50][143], dotarray[51][143], dotarray[52][143], dotarray[53][143], dotarray[54][143], dotarray[55][143], dotarray[56][143], dotarray[57][143], dotarray[58][143], dotarray[59][143], dotarray[60][143], dotarray[61][143], dotarray[62][143], dotarray[63][143], dotarray[64][143], dotarray[65][143], dotarray[66][143], dotarray[67][143], dotarray[68][143], dotarray[69][143], dotarray[70][143], dotarray[71][143], dotarray[72][143], dotarray[73][143], dotarray[74][143], dotarray[75][143], dotarray[76][143], dotarray[77][143], dotarray[78][143], dotarray[79][143], dotarray[80][143], dotarray[81][143], dotarray[82][143], dotarray[83][143], dotarray[84][143], dotarray[85][143], dotarray[86][143], dotarray[87][143], dotarray[88][143], dotarray[89][143], dotarray[90][143], dotarray[91][143], dotarray[92][143], dotarray[93][143], dotarray[94][143], dotarray[95][143], dotarray[96][143], dotarray[97][143], dotarray[98][143], dotarray[99][143], dotarray[100][143], dotarray[101][143], dotarray[102][143], dotarray[103][143], dotarray[104][143], dotarray[105][143], dotarray[106][143], dotarray[107][143], dotarray[108][143], dotarray[109][143], dotarray[110][143], dotarray[111][143], dotarray[112][143], dotarray[113][143], dotarray[114][143], dotarray[115][143], dotarray[116][143], dotarray[117][143], dotarray[118][143], dotarray[119][143], dotarray[120][143], dotarray[121][143], dotarray[122][143], dotarray[123][143], dotarray[124][143], dotarray[125][143], dotarray[126][143], dotarray[127][143]};
assign dot_col_144 = {dotarray[0][144], dotarray[1][144], dotarray[2][144], dotarray[3][144], dotarray[4][144], dotarray[5][144], dotarray[6][144], dotarray[7][144], dotarray[8][144], dotarray[9][144], dotarray[10][144], dotarray[11][144], dotarray[12][144], dotarray[13][144], dotarray[14][144], dotarray[15][144], dotarray[16][144], dotarray[17][144], dotarray[18][144], dotarray[19][144], dotarray[20][144], dotarray[21][144], dotarray[22][144], dotarray[23][144], dotarray[24][144], dotarray[25][144], dotarray[26][144], dotarray[27][144], dotarray[28][144], dotarray[29][144], dotarray[30][144], dotarray[31][144], dotarray[32][144], dotarray[33][144], dotarray[34][144], dotarray[35][144], dotarray[36][144], dotarray[37][144], dotarray[38][144], dotarray[39][144], dotarray[40][144], dotarray[41][144], dotarray[42][144], dotarray[43][144], dotarray[44][144], dotarray[45][144], dotarray[46][144], dotarray[47][144], dotarray[48][144], dotarray[49][144], dotarray[50][144], dotarray[51][144], dotarray[52][144], dotarray[53][144], dotarray[54][144], dotarray[55][144], dotarray[56][144], dotarray[57][144], dotarray[58][144], dotarray[59][144], dotarray[60][144], dotarray[61][144], dotarray[62][144], dotarray[63][144], dotarray[64][144], dotarray[65][144], dotarray[66][144], dotarray[67][144], dotarray[68][144], dotarray[69][144], dotarray[70][144], dotarray[71][144], dotarray[72][144], dotarray[73][144], dotarray[74][144], dotarray[75][144], dotarray[76][144], dotarray[77][144], dotarray[78][144], dotarray[79][144], dotarray[80][144], dotarray[81][144], dotarray[82][144], dotarray[83][144], dotarray[84][144], dotarray[85][144], dotarray[86][144], dotarray[87][144], dotarray[88][144], dotarray[89][144], dotarray[90][144], dotarray[91][144], dotarray[92][144], dotarray[93][144], dotarray[94][144], dotarray[95][144], dotarray[96][144], dotarray[97][144], dotarray[98][144], dotarray[99][144], dotarray[100][144], dotarray[101][144], dotarray[102][144], dotarray[103][144], dotarray[104][144], dotarray[105][144], dotarray[106][144], dotarray[107][144], dotarray[108][144], dotarray[109][144], dotarray[110][144], dotarray[111][144], dotarray[112][144], dotarray[113][144], dotarray[114][144], dotarray[115][144], dotarray[116][144], dotarray[117][144], dotarray[118][144], dotarray[119][144], dotarray[120][144], dotarray[121][144], dotarray[122][144], dotarray[123][144], dotarray[124][144], dotarray[125][144], dotarray[126][144], dotarray[127][144]};
assign dot_col_145 = {dotarray[0][145], dotarray[1][145], dotarray[2][145], dotarray[3][145], dotarray[4][145], dotarray[5][145], dotarray[6][145], dotarray[7][145], dotarray[8][145], dotarray[9][145], dotarray[10][145], dotarray[11][145], dotarray[12][145], dotarray[13][145], dotarray[14][145], dotarray[15][145], dotarray[16][145], dotarray[17][145], dotarray[18][145], dotarray[19][145], dotarray[20][145], dotarray[21][145], dotarray[22][145], dotarray[23][145], dotarray[24][145], dotarray[25][145], dotarray[26][145], dotarray[27][145], dotarray[28][145], dotarray[29][145], dotarray[30][145], dotarray[31][145], dotarray[32][145], dotarray[33][145], dotarray[34][145], dotarray[35][145], dotarray[36][145], dotarray[37][145], dotarray[38][145], dotarray[39][145], dotarray[40][145], dotarray[41][145], dotarray[42][145], dotarray[43][145], dotarray[44][145], dotarray[45][145], dotarray[46][145], dotarray[47][145], dotarray[48][145], dotarray[49][145], dotarray[50][145], dotarray[51][145], dotarray[52][145], dotarray[53][145], dotarray[54][145], dotarray[55][145], dotarray[56][145], dotarray[57][145], dotarray[58][145], dotarray[59][145], dotarray[60][145], dotarray[61][145], dotarray[62][145], dotarray[63][145], dotarray[64][145], dotarray[65][145], dotarray[66][145], dotarray[67][145], dotarray[68][145], dotarray[69][145], dotarray[70][145], dotarray[71][145], dotarray[72][145], dotarray[73][145], dotarray[74][145], dotarray[75][145], dotarray[76][145], dotarray[77][145], dotarray[78][145], dotarray[79][145], dotarray[80][145], dotarray[81][145], dotarray[82][145], dotarray[83][145], dotarray[84][145], dotarray[85][145], dotarray[86][145], dotarray[87][145], dotarray[88][145], dotarray[89][145], dotarray[90][145], dotarray[91][145], dotarray[92][145], dotarray[93][145], dotarray[94][145], dotarray[95][145], dotarray[96][145], dotarray[97][145], dotarray[98][145], dotarray[99][145], dotarray[100][145], dotarray[101][145], dotarray[102][145], dotarray[103][145], dotarray[104][145], dotarray[105][145], dotarray[106][145], dotarray[107][145], dotarray[108][145], dotarray[109][145], dotarray[110][145], dotarray[111][145], dotarray[112][145], dotarray[113][145], dotarray[114][145], dotarray[115][145], dotarray[116][145], dotarray[117][145], dotarray[118][145], dotarray[119][145], dotarray[120][145], dotarray[121][145], dotarray[122][145], dotarray[123][145], dotarray[124][145], dotarray[125][145], dotarray[126][145], dotarray[127][145]};
assign dot_col_146 = {dotarray[0][146], dotarray[1][146], dotarray[2][146], dotarray[3][146], dotarray[4][146], dotarray[5][146], dotarray[6][146], dotarray[7][146], dotarray[8][146], dotarray[9][146], dotarray[10][146], dotarray[11][146], dotarray[12][146], dotarray[13][146], dotarray[14][146], dotarray[15][146], dotarray[16][146], dotarray[17][146], dotarray[18][146], dotarray[19][146], dotarray[20][146], dotarray[21][146], dotarray[22][146], dotarray[23][146], dotarray[24][146], dotarray[25][146], dotarray[26][146], dotarray[27][146], dotarray[28][146], dotarray[29][146], dotarray[30][146], dotarray[31][146], dotarray[32][146], dotarray[33][146], dotarray[34][146], dotarray[35][146], dotarray[36][146], dotarray[37][146], dotarray[38][146], dotarray[39][146], dotarray[40][146], dotarray[41][146], dotarray[42][146], dotarray[43][146], dotarray[44][146], dotarray[45][146], dotarray[46][146], dotarray[47][146], dotarray[48][146], dotarray[49][146], dotarray[50][146], dotarray[51][146], dotarray[52][146], dotarray[53][146], dotarray[54][146], dotarray[55][146], dotarray[56][146], dotarray[57][146], dotarray[58][146], dotarray[59][146], dotarray[60][146], dotarray[61][146], dotarray[62][146], dotarray[63][146], dotarray[64][146], dotarray[65][146], dotarray[66][146], dotarray[67][146], dotarray[68][146], dotarray[69][146], dotarray[70][146], dotarray[71][146], dotarray[72][146], dotarray[73][146], dotarray[74][146], dotarray[75][146], dotarray[76][146], dotarray[77][146], dotarray[78][146], dotarray[79][146], dotarray[80][146], dotarray[81][146], dotarray[82][146], dotarray[83][146], dotarray[84][146], dotarray[85][146], dotarray[86][146], dotarray[87][146], dotarray[88][146], dotarray[89][146], dotarray[90][146], dotarray[91][146], dotarray[92][146], dotarray[93][146], dotarray[94][146], dotarray[95][146], dotarray[96][146], dotarray[97][146], dotarray[98][146], dotarray[99][146], dotarray[100][146], dotarray[101][146], dotarray[102][146], dotarray[103][146], dotarray[104][146], dotarray[105][146], dotarray[106][146], dotarray[107][146], dotarray[108][146], dotarray[109][146], dotarray[110][146], dotarray[111][146], dotarray[112][146], dotarray[113][146], dotarray[114][146], dotarray[115][146], dotarray[116][146], dotarray[117][146], dotarray[118][146], dotarray[119][146], dotarray[120][146], dotarray[121][146], dotarray[122][146], dotarray[123][146], dotarray[124][146], dotarray[125][146], dotarray[126][146], dotarray[127][146]};
assign dot_col_147 = {dotarray[0][147], dotarray[1][147], dotarray[2][147], dotarray[3][147], dotarray[4][147], dotarray[5][147], dotarray[6][147], dotarray[7][147], dotarray[8][147], dotarray[9][147], dotarray[10][147], dotarray[11][147], dotarray[12][147], dotarray[13][147], dotarray[14][147], dotarray[15][147], dotarray[16][147], dotarray[17][147], dotarray[18][147], dotarray[19][147], dotarray[20][147], dotarray[21][147], dotarray[22][147], dotarray[23][147], dotarray[24][147], dotarray[25][147], dotarray[26][147], dotarray[27][147], dotarray[28][147], dotarray[29][147], dotarray[30][147], dotarray[31][147], dotarray[32][147], dotarray[33][147], dotarray[34][147], dotarray[35][147], dotarray[36][147], dotarray[37][147], dotarray[38][147], dotarray[39][147], dotarray[40][147], dotarray[41][147], dotarray[42][147], dotarray[43][147], dotarray[44][147], dotarray[45][147], dotarray[46][147], dotarray[47][147], dotarray[48][147], dotarray[49][147], dotarray[50][147], dotarray[51][147], dotarray[52][147], dotarray[53][147], dotarray[54][147], dotarray[55][147], dotarray[56][147], dotarray[57][147], dotarray[58][147], dotarray[59][147], dotarray[60][147], dotarray[61][147], dotarray[62][147], dotarray[63][147], dotarray[64][147], dotarray[65][147], dotarray[66][147], dotarray[67][147], dotarray[68][147], dotarray[69][147], dotarray[70][147], dotarray[71][147], dotarray[72][147], dotarray[73][147], dotarray[74][147], dotarray[75][147], dotarray[76][147], dotarray[77][147], dotarray[78][147], dotarray[79][147], dotarray[80][147], dotarray[81][147], dotarray[82][147], dotarray[83][147], dotarray[84][147], dotarray[85][147], dotarray[86][147], dotarray[87][147], dotarray[88][147], dotarray[89][147], dotarray[90][147], dotarray[91][147], dotarray[92][147], dotarray[93][147], dotarray[94][147], dotarray[95][147], dotarray[96][147], dotarray[97][147], dotarray[98][147], dotarray[99][147], dotarray[100][147], dotarray[101][147], dotarray[102][147], dotarray[103][147], dotarray[104][147], dotarray[105][147], dotarray[106][147], dotarray[107][147], dotarray[108][147], dotarray[109][147], dotarray[110][147], dotarray[111][147], dotarray[112][147], dotarray[113][147], dotarray[114][147], dotarray[115][147], dotarray[116][147], dotarray[117][147], dotarray[118][147], dotarray[119][147], dotarray[120][147], dotarray[121][147], dotarray[122][147], dotarray[123][147], dotarray[124][147], dotarray[125][147], dotarray[126][147], dotarray[127][147]};
assign dot_col_148 = {dotarray[0][148], dotarray[1][148], dotarray[2][148], dotarray[3][148], dotarray[4][148], dotarray[5][148], dotarray[6][148], dotarray[7][148], dotarray[8][148], dotarray[9][148], dotarray[10][148], dotarray[11][148], dotarray[12][148], dotarray[13][148], dotarray[14][148], dotarray[15][148], dotarray[16][148], dotarray[17][148], dotarray[18][148], dotarray[19][148], dotarray[20][148], dotarray[21][148], dotarray[22][148], dotarray[23][148], dotarray[24][148], dotarray[25][148], dotarray[26][148], dotarray[27][148], dotarray[28][148], dotarray[29][148], dotarray[30][148], dotarray[31][148], dotarray[32][148], dotarray[33][148], dotarray[34][148], dotarray[35][148], dotarray[36][148], dotarray[37][148], dotarray[38][148], dotarray[39][148], dotarray[40][148], dotarray[41][148], dotarray[42][148], dotarray[43][148], dotarray[44][148], dotarray[45][148], dotarray[46][148], dotarray[47][148], dotarray[48][148], dotarray[49][148], dotarray[50][148], dotarray[51][148], dotarray[52][148], dotarray[53][148], dotarray[54][148], dotarray[55][148], dotarray[56][148], dotarray[57][148], dotarray[58][148], dotarray[59][148], dotarray[60][148], dotarray[61][148], dotarray[62][148], dotarray[63][148], dotarray[64][148], dotarray[65][148], dotarray[66][148], dotarray[67][148], dotarray[68][148], dotarray[69][148], dotarray[70][148], dotarray[71][148], dotarray[72][148], dotarray[73][148], dotarray[74][148], dotarray[75][148], dotarray[76][148], dotarray[77][148], dotarray[78][148], dotarray[79][148], dotarray[80][148], dotarray[81][148], dotarray[82][148], dotarray[83][148], dotarray[84][148], dotarray[85][148], dotarray[86][148], dotarray[87][148], dotarray[88][148], dotarray[89][148], dotarray[90][148], dotarray[91][148], dotarray[92][148], dotarray[93][148], dotarray[94][148], dotarray[95][148], dotarray[96][148], dotarray[97][148], dotarray[98][148], dotarray[99][148], dotarray[100][148], dotarray[101][148], dotarray[102][148], dotarray[103][148], dotarray[104][148], dotarray[105][148], dotarray[106][148], dotarray[107][148], dotarray[108][148], dotarray[109][148], dotarray[110][148], dotarray[111][148], dotarray[112][148], dotarray[113][148], dotarray[114][148], dotarray[115][148], dotarray[116][148], dotarray[117][148], dotarray[118][148], dotarray[119][148], dotarray[120][148], dotarray[121][148], dotarray[122][148], dotarray[123][148], dotarray[124][148], dotarray[125][148], dotarray[126][148], dotarray[127][148]};
assign dot_col_149 = {dotarray[0][149], dotarray[1][149], dotarray[2][149], dotarray[3][149], dotarray[4][149], dotarray[5][149], dotarray[6][149], dotarray[7][149], dotarray[8][149], dotarray[9][149], dotarray[10][149], dotarray[11][149], dotarray[12][149], dotarray[13][149], dotarray[14][149], dotarray[15][149], dotarray[16][149], dotarray[17][149], dotarray[18][149], dotarray[19][149], dotarray[20][149], dotarray[21][149], dotarray[22][149], dotarray[23][149], dotarray[24][149], dotarray[25][149], dotarray[26][149], dotarray[27][149], dotarray[28][149], dotarray[29][149], dotarray[30][149], dotarray[31][149], dotarray[32][149], dotarray[33][149], dotarray[34][149], dotarray[35][149], dotarray[36][149], dotarray[37][149], dotarray[38][149], dotarray[39][149], dotarray[40][149], dotarray[41][149], dotarray[42][149], dotarray[43][149], dotarray[44][149], dotarray[45][149], dotarray[46][149], dotarray[47][149], dotarray[48][149], dotarray[49][149], dotarray[50][149], dotarray[51][149], dotarray[52][149], dotarray[53][149], dotarray[54][149], dotarray[55][149], dotarray[56][149], dotarray[57][149], dotarray[58][149], dotarray[59][149], dotarray[60][149], dotarray[61][149], dotarray[62][149], dotarray[63][149], dotarray[64][149], dotarray[65][149], dotarray[66][149], dotarray[67][149], dotarray[68][149], dotarray[69][149], dotarray[70][149], dotarray[71][149], dotarray[72][149], dotarray[73][149], dotarray[74][149], dotarray[75][149], dotarray[76][149], dotarray[77][149], dotarray[78][149], dotarray[79][149], dotarray[80][149], dotarray[81][149], dotarray[82][149], dotarray[83][149], dotarray[84][149], dotarray[85][149], dotarray[86][149], dotarray[87][149], dotarray[88][149], dotarray[89][149], dotarray[90][149], dotarray[91][149], dotarray[92][149], dotarray[93][149], dotarray[94][149], dotarray[95][149], dotarray[96][149], dotarray[97][149], dotarray[98][149], dotarray[99][149], dotarray[100][149], dotarray[101][149], dotarray[102][149], dotarray[103][149], dotarray[104][149], dotarray[105][149], dotarray[106][149], dotarray[107][149], dotarray[108][149], dotarray[109][149], dotarray[110][149], dotarray[111][149], dotarray[112][149], dotarray[113][149], dotarray[114][149], dotarray[115][149], dotarray[116][149], dotarray[117][149], dotarray[118][149], dotarray[119][149], dotarray[120][149], dotarray[121][149], dotarray[122][149], dotarray[123][149], dotarray[124][149], dotarray[125][149], dotarray[126][149], dotarray[127][149]};
assign dot_col_150 = {dotarray[0][150], dotarray[1][150], dotarray[2][150], dotarray[3][150], dotarray[4][150], dotarray[5][150], dotarray[6][150], dotarray[7][150], dotarray[8][150], dotarray[9][150], dotarray[10][150], dotarray[11][150], dotarray[12][150], dotarray[13][150], dotarray[14][150], dotarray[15][150], dotarray[16][150], dotarray[17][150], dotarray[18][150], dotarray[19][150], dotarray[20][150], dotarray[21][150], dotarray[22][150], dotarray[23][150], dotarray[24][150], dotarray[25][150], dotarray[26][150], dotarray[27][150], dotarray[28][150], dotarray[29][150], dotarray[30][150], dotarray[31][150], dotarray[32][150], dotarray[33][150], dotarray[34][150], dotarray[35][150], dotarray[36][150], dotarray[37][150], dotarray[38][150], dotarray[39][150], dotarray[40][150], dotarray[41][150], dotarray[42][150], dotarray[43][150], dotarray[44][150], dotarray[45][150], dotarray[46][150], dotarray[47][150], dotarray[48][150], dotarray[49][150], dotarray[50][150], dotarray[51][150], dotarray[52][150], dotarray[53][150], dotarray[54][150], dotarray[55][150], dotarray[56][150], dotarray[57][150], dotarray[58][150], dotarray[59][150], dotarray[60][150], dotarray[61][150], dotarray[62][150], dotarray[63][150], dotarray[64][150], dotarray[65][150], dotarray[66][150], dotarray[67][150], dotarray[68][150], dotarray[69][150], dotarray[70][150], dotarray[71][150], dotarray[72][150], dotarray[73][150], dotarray[74][150], dotarray[75][150], dotarray[76][150], dotarray[77][150], dotarray[78][150], dotarray[79][150], dotarray[80][150], dotarray[81][150], dotarray[82][150], dotarray[83][150], dotarray[84][150], dotarray[85][150], dotarray[86][150], dotarray[87][150], dotarray[88][150], dotarray[89][150], dotarray[90][150], dotarray[91][150], dotarray[92][150], dotarray[93][150], dotarray[94][150], dotarray[95][150], dotarray[96][150], dotarray[97][150], dotarray[98][150], dotarray[99][150], dotarray[100][150], dotarray[101][150], dotarray[102][150], dotarray[103][150], dotarray[104][150], dotarray[105][150], dotarray[106][150], dotarray[107][150], dotarray[108][150], dotarray[109][150], dotarray[110][150], dotarray[111][150], dotarray[112][150], dotarray[113][150], dotarray[114][150], dotarray[115][150], dotarray[116][150], dotarray[117][150], dotarray[118][150], dotarray[119][150], dotarray[120][150], dotarray[121][150], dotarray[122][150], dotarray[123][150], dotarray[124][150], dotarray[125][150], dotarray[126][150], dotarray[127][150]};
assign dot_col_151 = {dotarray[0][151], dotarray[1][151], dotarray[2][151], dotarray[3][151], dotarray[4][151], dotarray[5][151], dotarray[6][151], dotarray[7][151], dotarray[8][151], dotarray[9][151], dotarray[10][151], dotarray[11][151], dotarray[12][151], dotarray[13][151], dotarray[14][151], dotarray[15][151], dotarray[16][151], dotarray[17][151], dotarray[18][151], dotarray[19][151], dotarray[20][151], dotarray[21][151], dotarray[22][151], dotarray[23][151], dotarray[24][151], dotarray[25][151], dotarray[26][151], dotarray[27][151], dotarray[28][151], dotarray[29][151], dotarray[30][151], dotarray[31][151], dotarray[32][151], dotarray[33][151], dotarray[34][151], dotarray[35][151], dotarray[36][151], dotarray[37][151], dotarray[38][151], dotarray[39][151], dotarray[40][151], dotarray[41][151], dotarray[42][151], dotarray[43][151], dotarray[44][151], dotarray[45][151], dotarray[46][151], dotarray[47][151], dotarray[48][151], dotarray[49][151], dotarray[50][151], dotarray[51][151], dotarray[52][151], dotarray[53][151], dotarray[54][151], dotarray[55][151], dotarray[56][151], dotarray[57][151], dotarray[58][151], dotarray[59][151], dotarray[60][151], dotarray[61][151], dotarray[62][151], dotarray[63][151], dotarray[64][151], dotarray[65][151], dotarray[66][151], dotarray[67][151], dotarray[68][151], dotarray[69][151], dotarray[70][151], dotarray[71][151], dotarray[72][151], dotarray[73][151], dotarray[74][151], dotarray[75][151], dotarray[76][151], dotarray[77][151], dotarray[78][151], dotarray[79][151], dotarray[80][151], dotarray[81][151], dotarray[82][151], dotarray[83][151], dotarray[84][151], dotarray[85][151], dotarray[86][151], dotarray[87][151], dotarray[88][151], dotarray[89][151], dotarray[90][151], dotarray[91][151], dotarray[92][151], dotarray[93][151], dotarray[94][151], dotarray[95][151], dotarray[96][151], dotarray[97][151], dotarray[98][151], dotarray[99][151], dotarray[100][151], dotarray[101][151], dotarray[102][151], dotarray[103][151], dotarray[104][151], dotarray[105][151], dotarray[106][151], dotarray[107][151], dotarray[108][151], dotarray[109][151], dotarray[110][151], dotarray[111][151], dotarray[112][151], dotarray[113][151], dotarray[114][151], dotarray[115][151], dotarray[116][151], dotarray[117][151], dotarray[118][151], dotarray[119][151], dotarray[120][151], dotarray[121][151], dotarray[122][151], dotarray[123][151], dotarray[124][151], dotarray[125][151], dotarray[126][151], dotarray[127][151]};
assign dot_col_152 = {dotarray[0][152], dotarray[1][152], dotarray[2][152], dotarray[3][152], dotarray[4][152], dotarray[5][152], dotarray[6][152], dotarray[7][152], dotarray[8][152], dotarray[9][152], dotarray[10][152], dotarray[11][152], dotarray[12][152], dotarray[13][152], dotarray[14][152], dotarray[15][152], dotarray[16][152], dotarray[17][152], dotarray[18][152], dotarray[19][152], dotarray[20][152], dotarray[21][152], dotarray[22][152], dotarray[23][152], dotarray[24][152], dotarray[25][152], dotarray[26][152], dotarray[27][152], dotarray[28][152], dotarray[29][152], dotarray[30][152], dotarray[31][152], dotarray[32][152], dotarray[33][152], dotarray[34][152], dotarray[35][152], dotarray[36][152], dotarray[37][152], dotarray[38][152], dotarray[39][152], dotarray[40][152], dotarray[41][152], dotarray[42][152], dotarray[43][152], dotarray[44][152], dotarray[45][152], dotarray[46][152], dotarray[47][152], dotarray[48][152], dotarray[49][152], dotarray[50][152], dotarray[51][152], dotarray[52][152], dotarray[53][152], dotarray[54][152], dotarray[55][152], dotarray[56][152], dotarray[57][152], dotarray[58][152], dotarray[59][152], dotarray[60][152], dotarray[61][152], dotarray[62][152], dotarray[63][152], dotarray[64][152], dotarray[65][152], dotarray[66][152], dotarray[67][152], dotarray[68][152], dotarray[69][152], dotarray[70][152], dotarray[71][152], dotarray[72][152], dotarray[73][152], dotarray[74][152], dotarray[75][152], dotarray[76][152], dotarray[77][152], dotarray[78][152], dotarray[79][152], dotarray[80][152], dotarray[81][152], dotarray[82][152], dotarray[83][152], dotarray[84][152], dotarray[85][152], dotarray[86][152], dotarray[87][152], dotarray[88][152], dotarray[89][152], dotarray[90][152], dotarray[91][152], dotarray[92][152], dotarray[93][152], dotarray[94][152], dotarray[95][152], dotarray[96][152], dotarray[97][152], dotarray[98][152], dotarray[99][152], dotarray[100][152], dotarray[101][152], dotarray[102][152], dotarray[103][152], dotarray[104][152], dotarray[105][152], dotarray[106][152], dotarray[107][152], dotarray[108][152], dotarray[109][152], dotarray[110][152], dotarray[111][152], dotarray[112][152], dotarray[113][152], dotarray[114][152], dotarray[115][152], dotarray[116][152], dotarray[117][152], dotarray[118][152], dotarray[119][152], dotarray[120][152], dotarray[121][152], dotarray[122][152], dotarray[123][152], dotarray[124][152], dotarray[125][152], dotarray[126][152], dotarray[127][152]};
assign dot_col_153 = {dotarray[0][153], dotarray[1][153], dotarray[2][153], dotarray[3][153], dotarray[4][153], dotarray[5][153], dotarray[6][153], dotarray[7][153], dotarray[8][153], dotarray[9][153], dotarray[10][153], dotarray[11][153], dotarray[12][153], dotarray[13][153], dotarray[14][153], dotarray[15][153], dotarray[16][153], dotarray[17][153], dotarray[18][153], dotarray[19][153], dotarray[20][153], dotarray[21][153], dotarray[22][153], dotarray[23][153], dotarray[24][153], dotarray[25][153], dotarray[26][153], dotarray[27][153], dotarray[28][153], dotarray[29][153], dotarray[30][153], dotarray[31][153], dotarray[32][153], dotarray[33][153], dotarray[34][153], dotarray[35][153], dotarray[36][153], dotarray[37][153], dotarray[38][153], dotarray[39][153], dotarray[40][153], dotarray[41][153], dotarray[42][153], dotarray[43][153], dotarray[44][153], dotarray[45][153], dotarray[46][153], dotarray[47][153], dotarray[48][153], dotarray[49][153], dotarray[50][153], dotarray[51][153], dotarray[52][153], dotarray[53][153], dotarray[54][153], dotarray[55][153], dotarray[56][153], dotarray[57][153], dotarray[58][153], dotarray[59][153], dotarray[60][153], dotarray[61][153], dotarray[62][153], dotarray[63][153], dotarray[64][153], dotarray[65][153], dotarray[66][153], dotarray[67][153], dotarray[68][153], dotarray[69][153], dotarray[70][153], dotarray[71][153], dotarray[72][153], dotarray[73][153], dotarray[74][153], dotarray[75][153], dotarray[76][153], dotarray[77][153], dotarray[78][153], dotarray[79][153], dotarray[80][153], dotarray[81][153], dotarray[82][153], dotarray[83][153], dotarray[84][153], dotarray[85][153], dotarray[86][153], dotarray[87][153], dotarray[88][153], dotarray[89][153], dotarray[90][153], dotarray[91][153], dotarray[92][153], dotarray[93][153], dotarray[94][153], dotarray[95][153], dotarray[96][153], dotarray[97][153], dotarray[98][153], dotarray[99][153], dotarray[100][153], dotarray[101][153], dotarray[102][153], dotarray[103][153], dotarray[104][153], dotarray[105][153], dotarray[106][153], dotarray[107][153], dotarray[108][153], dotarray[109][153], dotarray[110][153], dotarray[111][153], dotarray[112][153], dotarray[113][153], dotarray[114][153], dotarray[115][153], dotarray[116][153], dotarray[117][153], dotarray[118][153], dotarray[119][153], dotarray[120][153], dotarray[121][153], dotarray[122][153], dotarray[123][153], dotarray[124][153], dotarray[125][153], dotarray[126][153], dotarray[127][153]};
assign dot_col_154 = {dotarray[0][154], dotarray[1][154], dotarray[2][154], dotarray[3][154], dotarray[4][154], dotarray[5][154], dotarray[6][154], dotarray[7][154], dotarray[8][154], dotarray[9][154], dotarray[10][154], dotarray[11][154], dotarray[12][154], dotarray[13][154], dotarray[14][154], dotarray[15][154], dotarray[16][154], dotarray[17][154], dotarray[18][154], dotarray[19][154], dotarray[20][154], dotarray[21][154], dotarray[22][154], dotarray[23][154], dotarray[24][154], dotarray[25][154], dotarray[26][154], dotarray[27][154], dotarray[28][154], dotarray[29][154], dotarray[30][154], dotarray[31][154], dotarray[32][154], dotarray[33][154], dotarray[34][154], dotarray[35][154], dotarray[36][154], dotarray[37][154], dotarray[38][154], dotarray[39][154], dotarray[40][154], dotarray[41][154], dotarray[42][154], dotarray[43][154], dotarray[44][154], dotarray[45][154], dotarray[46][154], dotarray[47][154], dotarray[48][154], dotarray[49][154], dotarray[50][154], dotarray[51][154], dotarray[52][154], dotarray[53][154], dotarray[54][154], dotarray[55][154], dotarray[56][154], dotarray[57][154], dotarray[58][154], dotarray[59][154], dotarray[60][154], dotarray[61][154], dotarray[62][154], dotarray[63][154], dotarray[64][154], dotarray[65][154], dotarray[66][154], dotarray[67][154], dotarray[68][154], dotarray[69][154], dotarray[70][154], dotarray[71][154], dotarray[72][154], dotarray[73][154], dotarray[74][154], dotarray[75][154], dotarray[76][154], dotarray[77][154], dotarray[78][154], dotarray[79][154], dotarray[80][154], dotarray[81][154], dotarray[82][154], dotarray[83][154], dotarray[84][154], dotarray[85][154], dotarray[86][154], dotarray[87][154], dotarray[88][154], dotarray[89][154], dotarray[90][154], dotarray[91][154], dotarray[92][154], dotarray[93][154], dotarray[94][154], dotarray[95][154], dotarray[96][154], dotarray[97][154], dotarray[98][154], dotarray[99][154], dotarray[100][154], dotarray[101][154], dotarray[102][154], dotarray[103][154], dotarray[104][154], dotarray[105][154], dotarray[106][154], dotarray[107][154], dotarray[108][154], dotarray[109][154], dotarray[110][154], dotarray[111][154], dotarray[112][154], dotarray[113][154], dotarray[114][154], dotarray[115][154], dotarray[116][154], dotarray[117][154], dotarray[118][154], dotarray[119][154], dotarray[120][154], dotarray[121][154], dotarray[122][154], dotarray[123][154], dotarray[124][154], dotarray[125][154], dotarray[126][154], dotarray[127][154]};
assign dot_col_155 = {dotarray[0][155], dotarray[1][155], dotarray[2][155], dotarray[3][155], dotarray[4][155], dotarray[5][155], dotarray[6][155], dotarray[7][155], dotarray[8][155], dotarray[9][155], dotarray[10][155], dotarray[11][155], dotarray[12][155], dotarray[13][155], dotarray[14][155], dotarray[15][155], dotarray[16][155], dotarray[17][155], dotarray[18][155], dotarray[19][155], dotarray[20][155], dotarray[21][155], dotarray[22][155], dotarray[23][155], dotarray[24][155], dotarray[25][155], dotarray[26][155], dotarray[27][155], dotarray[28][155], dotarray[29][155], dotarray[30][155], dotarray[31][155], dotarray[32][155], dotarray[33][155], dotarray[34][155], dotarray[35][155], dotarray[36][155], dotarray[37][155], dotarray[38][155], dotarray[39][155], dotarray[40][155], dotarray[41][155], dotarray[42][155], dotarray[43][155], dotarray[44][155], dotarray[45][155], dotarray[46][155], dotarray[47][155], dotarray[48][155], dotarray[49][155], dotarray[50][155], dotarray[51][155], dotarray[52][155], dotarray[53][155], dotarray[54][155], dotarray[55][155], dotarray[56][155], dotarray[57][155], dotarray[58][155], dotarray[59][155], dotarray[60][155], dotarray[61][155], dotarray[62][155], dotarray[63][155], dotarray[64][155], dotarray[65][155], dotarray[66][155], dotarray[67][155], dotarray[68][155], dotarray[69][155], dotarray[70][155], dotarray[71][155], dotarray[72][155], dotarray[73][155], dotarray[74][155], dotarray[75][155], dotarray[76][155], dotarray[77][155], dotarray[78][155], dotarray[79][155], dotarray[80][155], dotarray[81][155], dotarray[82][155], dotarray[83][155], dotarray[84][155], dotarray[85][155], dotarray[86][155], dotarray[87][155], dotarray[88][155], dotarray[89][155], dotarray[90][155], dotarray[91][155], dotarray[92][155], dotarray[93][155], dotarray[94][155], dotarray[95][155], dotarray[96][155], dotarray[97][155], dotarray[98][155], dotarray[99][155], dotarray[100][155], dotarray[101][155], dotarray[102][155], dotarray[103][155], dotarray[104][155], dotarray[105][155], dotarray[106][155], dotarray[107][155], dotarray[108][155], dotarray[109][155], dotarray[110][155], dotarray[111][155], dotarray[112][155], dotarray[113][155], dotarray[114][155], dotarray[115][155], dotarray[116][155], dotarray[117][155], dotarray[118][155], dotarray[119][155], dotarray[120][155], dotarray[121][155], dotarray[122][155], dotarray[123][155], dotarray[124][155], dotarray[125][155], dotarray[126][155], dotarray[127][155]};
assign dot_col_156 = {dotarray[0][156], dotarray[1][156], dotarray[2][156], dotarray[3][156], dotarray[4][156], dotarray[5][156], dotarray[6][156], dotarray[7][156], dotarray[8][156], dotarray[9][156], dotarray[10][156], dotarray[11][156], dotarray[12][156], dotarray[13][156], dotarray[14][156], dotarray[15][156], dotarray[16][156], dotarray[17][156], dotarray[18][156], dotarray[19][156], dotarray[20][156], dotarray[21][156], dotarray[22][156], dotarray[23][156], dotarray[24][156], dotarray[25][156], dotarray[26][156], dotarray[27][156], dotarray[28][156], dotarray[29][156], dotarray[30][156], dotarray[31][156], dotarray[32][156], dotarray[33][156], dotarray[34][156], dotarray[35][156], dotarray[36][156], dotarray[37][156], dotarray[38][156], dotarray[39][156], dotarray[40][156], dotarray[41][156], dotarray[42][156], dotarray[43][156], dotarray[44][156], dotarray[45][156], dotarray[46][156], dotarray[47][156], dotarray[48][156], dotarray[49][156], dotarray[50][156], dotarray[51][156], dotarray[52][156], dotarray[53][156], dotarray[54][156], dotarray[55][156], dotarray[56][156], dotarray[57][156], dotarray[58][156], dotarray[59][156], dotarray[60][156], dotarray[61][156], dotarray[62][156], dotarray[63][156], dotarray[64][156], dotarray[65][156], dotarray[66][156], dotarray[67][156], dotarray[68][156], dotarray[69][156], dotarray[70][156], dotarray[71][156], dotarray[72][156], dotarray[73][156], dotarray[74][156], dotarray[75][156], dotarray[76][156], dotarray[77][156], dotarray[78][156], dotarray[79][156], dotarray[80][156], dotarray[81][156], dotarray[82][156], dotarray[83][156], dotarray[84][156], dotarray[85][156], dotarray[86][156], dotarray[87][156], dotarray[88][156], dotarray[89][156], dotarray[90][156], dotarray[91][156], dotarray[92][156], dotarray[93][156], dotarray[94][156], dotarray[95][156], dotarray[96][156], dotarray[97][156], dotarray[98][156], dotarray[99][156], dotarray[100][156], dotarray[101][156], dotarray[102][156], dotarray[103][156], dotarray[104][156], dotarray[105][156], dotarray[106][156], dotarray[107][156], dotarray[108][156], dotarray[109][156], dotarray[110][156], dotarray[111][156], dotarray[112][156], dotarray[113][156], dotarray[114][156], dotarray[115][156], dotarray[116][156], dotarray[117][156], dotarray[118][156], dotarray[119][156], dotarray[120][156], dotarray[121][156], dotarray[122][156], dotarray[123][156], dotarray[124][156], dotarray[125][156], dotarray[126][156], dotarray[127][156]};
assign dot_col_157 = {dotarray[0][157], dotarray[1][157], dotarray[2][157], dotarray[3][157], dotarray[4][157], dotarray[5][157], dotarray[6][157], dotarray[7][157], dotarray[8][157], dotarray[9][157], dotarray[10][157], dotarray[11][157], dotarray[12][157], dotarray[13][157], dotarray[14][157], dotarray[15][157], dotarray[16][157], dotarray[17][157], dotarray[18][157], dotarray[19][157], dotarray[20][157], dotarray[21][157], dotarray[22][157], dotarray[23][157], dotarray[24][157], dotarray[25][157], dotarray[26][157], dotarray[27][157], dotarray[28][157], dotarray[29][157], dotarray[30][157], dotarray[31][157], dotarray[32][157], dotarray[33][157], dotarray[34][157], dotarray[35][157], dotarray[36][157], dotarray[37][157], dotarray[38][157], dotarray[39][157], dotarray[40][157], dotarray[41][157], dotarray[42][157], dotarray[43][157], dotarray[44][157], dotarray[45][157], dotarray[46][157], dotarray[47][157], dotarray[48][157], dotarray[49][157], dotarray[50][157], dotarray[51][157], dotarray[52][157], dotarray[53][157], dotarray[54][157], dotarray[55][157], dotarray[56][157], dotarray[57][157], dotarray[58][157], dotarray[59][157], dotarray[60][157], dotarray[61][157], dotarray[62][157], dotarray[63][157], dotarray[64][157], dotarray[65][157], dotarray[66][157], dotarray[67][157], dotarray[68][157], dotarray[69][157], dotarray[70][157], dotarray[71][157], dotarray[72][157], dotarray[73][157], dotarray[74][157], dotarray[75][157], dotarray[76][157], dotarray[77][157], dotarray[78][157], dotarray[79][157], dotarray[80][157], dotarray[81][157], dotarray[82][157], dotarray[83][157], dotarray[84][157], dotarray[85][157], dotarray[86][157], dotarray[87][157], dotarray[88][157], dotarray[89][157], dotarray[90][157], dotarray[91][157], dotarray[92][157], dotarray[93][157], dotarray[94][157], dotarray[95][157], dotarray[96][157], dotarray[97][157], dotarray[98][157], dotarray[99][157], dotarray[100][157], dotarray[101][157], dotarray[102][157], dotarray[103][157], dotarray[104][157], dotarray[105][157], dotarray[106][157], dotarray[107][157], dotarray[108][157], dotarray[109][157], dotarray[110][157], dotarray[111][157], dotarray[112][157], dotarray[113][157], dotarray[114][157], dotarray[115][157], dotarray[116][157], dotarray[117][157], dotarray[118][157], dotarray[119][157], dotarray[120][157], dotarray[121][157], dotarray[122][157], dotarray[123][157], dotarray[124][157], dotarray[125][157], dotarray[126][157], dotarray[127][157]};
assign dot_col_158 = {dotarray[0][158], dotarray[1][158], dotarray[2][158], dotarray[3][158], dotarray[4][158], dotarray[5][158], dotarray[6][158], dotarray[7][158], dotarray[8][158], dotarray[9][158], dotarray[10][158], dotarray[11][158], dotarray[12][158], dotarray[13][158], dotarray[14][158], dotarray[15][158], dotarray[16][158], dotarray[17][158], dotarray[18][158], dotarray[19][158], dotarray[20][158], dotarray[21][158], dotarray[22][158], dotarray[23][158], dotarray[24][158], dotarray[25][158], dotarray[26][158], dotarray[27][158], dotarray[28][158], dotarray[29][158], dotarray[30][158], dotarray[31][158], dotarray[32][158], dotarray[33][158], dotarray[34][158], dotarray[35][158], dotarray[36][158], dotarray[37][158], dotarray[38][158], dotarray[39][158], dotarray[40][158], dotarray[41][158], dotarray[42][158], dotarray[43][158], dotarray[44][158], dotarray[45][158], dotarray[46][158], dotarray[47][158], dotarray[48][158], dotarray[49][158], dotarray[50][158], dotarray[51][158], dotarray[52][158], dotarray[53][158], dotarray[54][158], dotarray[55][158], dotarray[56][158], dotarray[57][158], dotarray[58][158], dotarray[59][158], dotarray[60][158], dotarray[61][158], dotarray[62][158], dotarray[63][158], dotarray[64][158], dotarray[65][158], dotarray[66][158], dotarray[67][158], dotarray[68][158], dotarray[69][158], dotarray[70][158], dotarray[71][158], dotarray[72][158], dotarray[73][158], dotarray[74][158], dotarray[75][158], dotarray[76][158], dotarray[77][158], dotarray[78][158], dotarray[79][158], dotarray[80][158], dotarray[81][158], dotarray[82][158], dotarray[83][158], dotarray[84][158], dotarray[85][158], dotarray[86][158], dotarray[87][158], dotarray[88][158], dotarray[89][158], dotarray[90][158], dotarray[91][158], dotarray[92][158], dotarray[93][158], dotarray[94][158], dotarray[95][158], dotarray[96][158], dotarray[97][158], dotarray[98][158], dotarray[99][158], dotarray[100][158], dotarray[101][158], dotarray[102][158], dotarray[103][158], dotarray[104][158], dotarray[105][158], dotarray[106][158], dotarray[107][158], dotarray[108][158], dotarray[109][158], dotarray[110][158], dotarray[111][158], dotarray[112][158], dotarray[113][158], dotarray[114][158], dotarray[115][158], dotarray[116][158], dotarray[117][158], dotarray[118][158], dotarray[119][158], dotarray[120][158], dotarray[121][158], dotarray[122][158], dotarray[123][158], dotarray[124][158], dotarray[125][158], dotarray[126][158], dotarray[127][158]};
assign dot_col_159 = {dotarray[0][159], dotarray[1][159], dotarray[2][159], dotarray[3][159], dotarray[4][159], dotarray[5][159], dotarray[6][159], dotarray[7][159], dotarray[8][159], dotarray[9][159], dotarray[10][159], dotarray[11][159], dotarray[12][159], dotarray[13][159], dotarray[14][159], dotarray[15][159], dotarray[16][159], dotarray[17][159], dotarray[18][159], dotarray[19][159], dotarray[20][159], dotarray[21][159], dotarray[22][159], dotarray[23][159], dotarray[24][159], dotarray[25][159], dotarray[26][159], dotarray[27][159], dotarray[28][159], dotarray[29][159], dotarray[30][159], dotarray[31][159], dotarray[32][159], dotarray[33][159], dotarray[34][159], dotarray[35][159], dotarray[36][159], dotarray[37][159], dotarray[38][159], dotarray[39][159], dotarray[40][159], dotarray[41][159], dotarray[42][159], dotarray[43][159], dotarray[44][159], dotarray[45][159], dotarray[46][159], dotarray[47][159], dotarray[48][159], dotarray[49][159], dotarray[50][159], dotarray[51][159], dotarray[52][159], dotarray[53][159], dotarray[54][159], dotarray[55][159], dotarray[56][159], dotarray[57][159], dotarray[58][159], dotarray[59][159], dotarray[60][159], dotarray[61][159], dotarray[62][159], dotarray[63][159], dotarray[64][159], dotarray[65][159], dotarray[66][159], dotarray[67][159], dotarray[68][159], dotarray[69][159], dotarray[70][159], dotarray[71][159], dotarray[72][159], dotarray[73][159], dotarray[74][159], dotarray[75][159], dotarray[76][159], dotarray[77][159], dotarray[78][159], dotarray[79][159], dotarray[80][159], dotarray[81][159], dotarray[82][159], dotarray[83][159], dotarray[84][159], dotarray[85][159], dotarray[86][159], dotarray[87][159], dotarray[88][159], dotarray[89][159], dotarray[90][159], dotarray[91][159], dotarray[92][159], dotarray[93][159], dotarray[94][159], dotarray[95][159], dotarray[96][159], dotarray[97][159], dotarray[98][159], dotarray[99][159], dotarray[100][159], dotarray[101][159], dotarray[102][159], dotarray[103][159], dotarray[104][159], dotarray[105][159], dotarray[106][159], dotarray[107][159], dotarray[108][159], dotarray[109][159], dotarray[110][159], dotarray[111][159], dotarray[112][159], dotarray[113][159], dotarray[114][159], dotarray[115][159], dotarray[116][159], dotarray[117][159], dotarray[118][159], dotarray[119][159], dotarray[120][159], dotarray[121][159], dotarray[122][159], dotarray[123][159], dotarray[124][159], dotarray[125][159], dotarray[126][159], dotarray[127][159]};
assign dot_col_160 = {dotarray[0][160], dotarray[1][160], dotarray[2][160], dotarray[3][160], dotarray[4][160], dotarray[5][160], dotarray[6][160], dotarray[7][160], dotarray[8][160], dotarray[9][160], dotarray[10][160], dotarray[11][160], dotarray[12][160], dotarray[13][160], dotarray[14][160], dotarray[15][160], dotarray[16][160], dotarray[17][160], dotarray[18][160], dotarray[19][160], dotarray[20][160], dotarray[21][160], dotarray[22][160], dotarray[23][160], dotarray[24][160], dotarray[25][160], dotarray[26][160], dotarray[27][160], dotarray[28][160], dotarray[29][160], dotarray[30][160], dotarray[31][160], dotarray[32][160], dotarray[33][160], dotarray[34][160], dotarray[35][160], dotarray[36][160], dotarray[37][160], dotarray[38][160], dotarray[39][160], dotarray[40][160], dotarray[41][160], dotarray[42][160], dotarray[43][160], dotarray[44][160], dotarray[45][160], dotarray[46][160], dotarray[47][160], dotarray[48][160], dotarray[49][160], dotarray[50][160], dotarray[51][160], dotarray[52][160], dotarray[53][160], dotarray[54][160], dotarray[55][160], dotarray[56][160], dotarray[57][160], dotarray[58][160], dotarray[59][160], dotarray[60][160], dotarray[61][160], dotarray[62][160], dotarray[63][160], dotarray[64][160], dotarray[65][160], dotarray[66][160], dotarray[67][160], dotarray[68][160], dotarray[69][160], dotarray[70][160], dotarray[71][160], dotarray[72][160], dotarray[73][160], dotarray[74][160], dotarray[75][160], dotarray[76][160], dotarray[77][160], dotarray[78][160], dotarray[79][160], dotarray[80][160], dotarray[81][160], dotarray[82][160], dotarray[83][160], dotarray[84][160], dotarray[85][160], dotarray[86][160], dotarray[87][160], dotarray[88][160], dotarray[89][160], dotarray[90][160], dotarray[91][160], dotarray[92][160], dotarray[93][160], dotarray[94][160], dotarray[95][160], dotarray[96][160], dotarray[97][160], dotarray[98][160], dotarray[99][160], dotarray[100][160], dotarray[101][160], dotarray[102][160], dotarray[103][160], dotarray[104][160], dotarray[105][160], dotarray[106][160], dotarray[107][160], dotarray[108][160], dotarray[109][160], dotarray[110][160], dotarray[111][160], dotarray[112][160], dotarray[113][160], dotarray[114][160], dotarray[115][160], dotarray[116][160], dotarray[117][160], dotarray[118][160], dotarray[119][160], dotarray[120][160], dotarray[121][160], dotarray[122][160], dotarray[123][160], dotarray[124][160], dotarray[125][160], dotarray[126][160], dotarray[127][160]};
assign dot_col_161 = {dotarray[0][161], dotarray[1][161], dotarray[2][161], dotarray[3][161], dotarray[4][161], dotarray[5][161], dotarray[6][161], dotarray[7][161], dotarray[8][161], dotarray[9][161], dotarray[10][161], dotarray[11][161], dotarray[12][161], dotarray[13][161], dotarray[14][161], dotarray[15][161], dotarray[16][161], dotarray[17][161], dotarray[18][161], dotarray[19][161], dotarray[20][161], dotarray[21][161], dotarray[22][161], dotarray[23][161], dotarray[24][161], dotarray[25][161], dotarray[26][161], dotarray[27][161], dotarray[28][161], dotarray[29][161], dotarray[30][161], dotarray[31][161], dotarray[32][161], dotarray[33][161], dotarray[34][161], dotarray[35][161], dotarray[36][161], dotarray[37][161], dotarray[38][161], dotarray[39][161], dotarray[40][161], dotarray[41][161], dotarray[42][161], dotarray[43][161], dotarray[44][161], dotarray[45][161], dotarray[46][161], dotarray[47][161], dotarray[48][161], dotarray[49][161], dotarray[50][161], dotarray[51][161], dotarray[52][161], dotarray[53][161], dotarray[54][161], dotarray[55][161], dotarray[56][161], dotarray[57][161], dotarray[58][161], dotarray[59][161], dotarray[60][161], dotarray[61][161], dotarray[62][161], dotarray[63][161], dotarray[64][161], dotarray[65][161], dotarray[66][161], dotarray[67][161], dotarray[68][161], dotarray[69][161], dotarray[70][161], dotarray[71][161], dotarray[72][161], dotarray[73][161], dotarray[74][161], dotarray[75][161], dotarray[76][161], dotarray[77][161], dotarray[78][161], dotarray[79][161], dotarray[80][161], dotarray[81][161], dotarray[82][161], dotarray[83][161], dotarray[84][161], dotarray[85][161], dotarray[86][161], dotarray[87][161], dotarray[88][161], dotarray[89][161], dotarray[90][161], dotarray[91][161], dotarray[92][161], dotarray[93][161], dotarray[94][161], dotarray[95][161], dotarray[96][161], dotarray[97][161], dotarray[98][161], dotarray[99][161], dotarray[100][161], dotarray[101][161], dotarray[102][161], dotarray[103][161], dotarray[104][161], dotarray[105][161], dotarray[106][161], dotarray[107][161], dotarray[108][161], dotarray[109][161], dotarray[110][161], dotarray[111][161], dotarray[112][161], dotarray[113][161], dotarray[114][161], dotarray[115][161], dotarray[116][161], dotarray[117][161], dotarray[118][161], dotarray[119][161], dotarray[120][161], dotarray[121][161], dotarray[122][161], dotarray[123][161], dotarray[124][161], dotarray[125][161], dotarray[126][161], dotarray[127][161]};
assign dot_col_162 = {dotarray[0][162], dotarray[1][162], dotarray[2][162], dotarray[3][162], dotarray[4][162], dotarray[5][162], dotarray[6][162], dotarray[7][162], dotarray[8][162], dotarray[9][162], dotarray[10][162], dotarray[11][162], dotarray[12][162], dotarray[13][162], dotarray[14][162], dotarray[15][162], dotarray[16][162], dotarray[17][162], dotarray[18][162], dotarray[19][162], dotarray[20][162], dotarray[21][162], dotarray[22][162], dotarray[23][162], dotarray[24][162], dotarray[25][162], dotarray[26][162], dotarray[27][162], dotarray[28][162], dotarray[29][162], dotarray[30][162], dotarray[31][162], dotarray[32][162], dotarray[33][162], dotarray[34][162], dotarray[35][162], dotarray[36][162], dotarray[37][162], dotarray[38][162], dotarray[39][162], dotarray[40][162], dotarray[41][162], dotarray[42][162], dotarray[43][162], dotarray[44][162], dotarray[45][162], dotarray[46][162], dotarray[47][162], dotarray[48][162], dotarray[49][162], dotarray[50][162], dotarray[51][162], dotarray[52][162], dotarray[53][162], dotarray[54][162], dotarray[55][162], dotarray[56][162], dotarray[57][162], dotarray[58][162], dotarray[59][162], dotarray[60][162], dotarray[61][162], dotarray[62][162], dotarray[63][162], dotarray[64][162], dotarray[65][162], dotarray[66][162], dotarray[67][162], dotarray[68][162], dotarray[69][162], dotarray[70][162], dotarray[71][162], dotarray[72][162], dotarray[73][162], dotarray[74][162], dotarray[75][162], dotarray[76][162], dotarray[77][162], dotarray[78][162], dotarray[79][162], dotarray[80][162], dotarray[81][162], dotarray[82][162], dotarray[83][162], dotarray[84][162], dotarray[85][162], dotarray[86][162], dotarray[87][162], dotarray[88][162], dotarray[89][162], dotarray[90][162], dotarray[91][162], dotarray[92][162], dotarray[93][162], dotarray[94][162], dotarray[95][162], dotarray[96][162], dotarray[97][162], dotarray[98][162], dotarray[99][162], dotarray[100][162], dotarray[101][162], dotarray[102][162], dotarray[103][162], dotarray[104][162], dotarray[105][162], dotarray[106][162], dotarray[107][162], dotarray[108][162], dotarray[109][162], dotarray[110][162], dotarray[111][162], dotarray[112][162], dotarray[113][162], dotarray[114][162], dotarray[115][162], dotarray[116][162], dotarray[117][162], dotarray[118][162], dotarray[119][162], dotarray[120][162], dotarray[121][162], dotarray[122][162], dotarray[123][162], dotarray[124][162], dotarray[125][162], dotarray[126][162], dotarray[127][162]};
assign dot_col_163 = {dotarray[0][163], dotarray[1][163], dotarray[2][163], dotarray[3][163], dotarray[4][163], dotarray[5][163], dotarray[6][163], dotarray[7][163], dotarray[8][163], dotarray[9][163], dotarray[10][163], dotarray[11][163], dotarray[12][163], dotarray[13][163], dotarray[14][163], dotarray[15][163], dotarray[16][163], dotarray[17][163], dotarray[18][163], dotarray[19][163], dotarray[20][163], dotarray[21][163], dotarray[22][163], dotarray[23][163], dotarray[24][163], dotarray[25][163], dotarray[26][163], dotarray[27][163], dotarray[28][163], dotarray[29][163], dotarray[30][163], dotarray[31][163], dotarray[32][163], dotarray[33][163], dotarray[34][163], dotarray[35][163], dotarray[36][163], dotarray[37][163], dotarray[38][163], dotarray[39][163], dotarray[40][163], dotarray[41][163], dotarray[42][163], dotarray[43][163], dotarray[44][163], dotarray[45][163], dotarray[46][163], dotarray[47][163], dotarray[48][163], dotarray[49][163], dotarray[50][163], dotarray[51][163], dotarray[52][163], dotarray[53][163], dotarray[54][163], dotarray[55][163], dotarray[56][163], dotarray[57][163], dotarray[58][163], dotarray[59][163], dotarray[60][163], dotarray[61][163], dotarray[62][163], dotarray[63][163], dotarray[64][163], dotarray[65][163], dotarray[66][163], dotarray[67][163], dotarray[68][163], dotarray[69][163], dotarray[70][163], dotarray[71][163], dotarray[72][163], dotarray[73][163], dotarray[74][163], dotarray[75][163], dotarray[76][163], dotarray[77][163], dotarray[78][163], dotarray[79][163], dotarray[80][163], dotarray[81][163], dotarray[82][163], dotarray[83][163], dotarray[84][163], dotarray[85][163], dotarray[86][163], dotarray[87][163], dotarray[88][163], dotarray[89][163], dotarray[90][163], dotarray[91][163], dotarray[92][163], dotarray[93][163], dotarray[94][163], dotarray[95][163], dotarray[96][163], dotarray[97][163], dotarray[98][163], dotarray[99][163], dotarray[100][163], dotarray[101][163], dotarray[102][163], dotarray[103][163], dotarray[104][163], dotarray[105][163], dotarray[106][163], dotarray[107][163], dotarray[108][163], dotarray[109][163], dotarray[110][163], dotarray[111][163], dotarray[112][163], dotarray[113][163], dotarray[114][163], dotarray[115][163], dotarray[116][163], dotarray[117][163], dotarray[118][163], dotarray[119][163], dotarray[120][163], dotarray[121][163], dotarray[122][163], dotarray[123][163], dotarray[124][163], dotarray[125][163], dotarray[126][163], dotarray[127][163]};
assign dot_col_164 = {dotarray[0][164], dotarray[1][164], dotarray[2][164], dotarray[3][164], dotarray[4][164], dotarray[5][164], dotarray[6][164], dotarray[7][164], dotarray[8][164], dotarray[9][164], dotarray[10][164], dotarray[11][164], dotarray[12][164], dotarray[13][164], dotarray[14][164], dotarray[15][164], dotarray[16][164], dotarray[17][164], dotarray[18][164], dotarray[19][164], dotarray[20][164], dotarray[21][164], dotarray[22][164], dotarray[23][164], dotarray[24][164], dotarray[25][164], dotarray[26][164], dotarray[27][164], dotarray[28][164], dotarray[29][164], dotarray[30][164], dotarray[31][164], dotarray[32][164], dotarray[33][164], dotarray[34][164], dotarray[35][164], dotarray[36][164], dotarray[37][164], dotarray[38][164], dotarray[39][164], dotarray[40][164], dotarray[41][164], dotarray[42][164], dotarray[43][164], dotarray[44][164], dotarray[45][164], dotarray[46][164], dotarray[47][164], dotarray[48][164], dotarray[49][164], dotarray[50][164], dotarray[51][164], dotarray[52][164], dotarray[53][164], dotarray[54][164], dotarray[55][164], dotarray[56][164], dotarray[57][164], dotarray[58][164], dotarray[59][164], dotarray[60][164], dotarray[61][164], dotarray[62][164], dotarray[63][164], dotarray[64][164], dotarray[65][164], dotarray[66][164], dotarray[67][164], dotarray[68][164], dotarray[69][164], dotarray[70][164], dotarray[71][164], dotarray[72][164], dotarray[73][164], dotarray[74][164], dotarray[75][164], dotarray[76][164], dotarray[77][164], dotarray[78][164], dotarray[79][164], dotarray[80][164], dotarray[81][164], dotarray[82][164], dotarray[83][164], dotarray[84][164], dotarray[85][164], dotarray[86][164], dotarray[87][164], dotarray[88][164], dotarray[89][164], dotarray[90][164], dotarray[91][164], dotarray[92][164], dotarray[93][164], dotarray[94][164], dotarray[95][164], dotarray[96][164], dotarray[97][164], dotarray[98][164], dotarray[99][164], dotarray[100][164], dotarray[101][164], dotarray[102][164], dotarray[103][164], dotarray[104][164], dotarray[105][164], dotarray[106][164], dotarray[107][164], dotarray[108][164], dotarray[109][164], dotarray[110][164], dotarray[111][164], dotarray[112][164], dotarray[113][164], dotarray[114][164], dotarray[115][164], dotarray[116][164], dotarray[117][164], dotarray[118][164], dotarray[119][164], dotarray[120][164], dotarray[121][164], dotarray[122][164], dotarray[123][164], dotarray[124][164], dotarray[125][164], dotarray[126][164], dotarray[127][164]};
assign dot_col_165 = {dotarray[0][165], dotarray[1][165], dotarray[2][165], dotarray[3][165], dotarray[4][165], dotarray[5][165], dotarray[6][165], dotarray[7][165], dotarray[8][165], dotarray[9][165], dotarray[10][165], dotarray[11][165], dotarray[12][165], dotarray[13][165], dotarray[14][165], dotarray[15][165], dotarray[16][165], dotarray[17][165], dotarray[18][165], dotarray[19][165], dotarray[20][165], dotarray[21][165], dotarray[22][165], dotarray[23][165], dotarray[24][165], dotarray[25][165], dotarray[26][165], dotarray[27][165], dotarray[28][165], dotarray[29][165], dotarray[30][165], dotarray[31][165], dotarray[32][165], dotarray[33][165], dotarray[34][165], dotarray[35][165], dotarray[36][165], dotarray[37][165], dotarray[38][165], dotarray[39][165], dotarray[40][165], dotarray[41][165], dotarray[42][165], dotarray[43][165], dotarray[44][165], dotarray[45][165], dotarray[46][165], dotarray[47][165], dotarray[48][165], dotarray[49][165], dotarray[50][165], dotarray[51][165], dotarray[52][165], dotarray[53][165], dotarray[54][165], dotarray[55][165], dotarray[56][165], dotarray[57][165], dotarray[58][165], dotarray[59][165], dotarray[60][165], dotarray[61][165], dotarray[62][165], dotarray[63][165], dotarray[64][165], dotarray[65][165], dotarray[66][165], dotarray[67][165], dotarray[68][165], dotarray[69][165], dotarray[70][165], dotarray[71][165], dotarray[72][165], dotarray[73][165], dotarray[74][165], dotarray[75][165], dotarray[76][165], dotarray[77][165], dotarray[78][165], dotarray[79][165], dotarray[80][165], dotarray[81][165], dotarray[82][165], dotarray[83][165], dotarray[84][165], dotarray[85][165], dotarray[86][165], dotarray[87][165], dotarray[88][165], dotarray[89][165], dotarray[90][165], dotarray[91][165], dotarray[92][165], dotarray[93][165], dotarray[94][165], dotarray[95][165], dotarray[96][165], dotarray[97][165], dotarray[98][165], dotarray[99][165], dotarray[100][165], dotarray[101][165], dotarray[102][165], dotarray[103][165], dotarray[104][165], dotarray[105][165], dotarray[106][165], dotarray[107][165], dotarray[108][165], dotarray[109][165], dotarray[110][165], dotarray[111][165], dotarray[112][165], dotarray[113][165], dotarray[114][165], dotarray[115][165], dotarray[116][165], dotarray[117][165], dotarray[118][165], dotarray[119][165], dotarray[120][165], dotarray[121][165], dotarray[122][165], dotarray[123][165], dotarray[124][165], dotarray[125][165], dotarray[126][165], dotarray[127][165]};
assign dot_col_166 = {dotarray[0][166], dotarray[1][166], dotarray[2][166], dotarray[3][166], dotarray[4][166], dotarray[5][166], dotarray[6][166], dotarray[7][166], dotarray[8][166], dotarray[9][166], dotarray[10][166], dotarray[11][166], dotarray[12][166], dotarray[13][166], dotarray[14][166], dotarray[15][166], dotarray[16][166], dotarray[17][166], dotarray[18][166], dotarray[19][166], dotarray[20][166], dotarray[21][166], dotarray[22][166], dotarray[23][166], dotarray[24][166], dotarray[25][166], dotarray[26][166], dotarray[27][166], dotarray[28][166], dotarray[29][166], dotarray[30][166], dotarray[31][166], dotarray[32][166], dotarray[33][166], dotarray[34][166], dotarray[35][166], dotarray[36][166], dotarray[37][166], dotarray[38][166], dotarray[39][166], dotarray[40][166], dotarray[41][166], dotarray[42][166], dotarray[43][166], dotarray[44][166], dotarray[45][166], dotarray[46][166], dotarray[47][166], dotarray[48][166], dotarray[49][166], dotarray[50][166], dotarray[51][166], dotarray[52][166], dotarray[53][166], dotarray[54][166], dotarray[55][166], dotarray[56][166], dotarray[57][166], dotarray[58][166], dotarray[59][166], dotarray[60][166], dotarray[61][166], dotarray[62][166], dotarray[63][166], dotarray[64][166], dotarray[65][166], dotarray[66][166], dotarray[67][166], dotarray[68][166], dotarray[69][166], dotarray[70][166], dotarray[71][166], dotarray[72][166], dotarray[73][166], dotarray[74][166], dotarray[75][166], dotarray[76][166], dotarray[77][166], dotarray[78][166], dotarray[79][166], dotarray[80][166], dotarray[81][166], dotarray[82][166], dotarray[83][166], dotarray[84][166], dotarray[85][166], dotarray[86][166], dotarray[87][166], dotarray[88][166], dotarray[89][166], dotarray[90][166], dotarray[91][166], dotarray[92][166], dotarray[93][166], dotarray[94][166], dotarray[95][166], dotarray[96][166], dotarray[97][166], dotarray[98][166], dotarray[99][166], dotarray[100][166], dotarray[101][166], dotarray[102][166], dotarray[103][166], dotarray[104][166], dotarray[105][166], dotarray[106][166], dotarray[107][166], dotarray[108][166], dotarray[109][166], dotarray[110][166], dotarray[111][166], dotarray[112][166], dotarray[113][166], dotarray[114][166], dotarray[115][166], dotarray[116][166], dotarray[117][166], dotarray[118][166], dotarray[119][166], dotarray[120][166], dotarray[121][166], dotarray[122][166], dotarray[123][166], dotarray[124][166], dotarray[125][166], dotarray[126][166], dotarray[127][166]};
assign dot_col_167 = {dotarray[0][167], dotarray[1][167], dotarray[2][167], dotarray[3][167], dotarray[4][167], dotarray[5][167], dotarray[6][167], dotarray[7][167], dotarray[8][167], dotarray[9][167], dotarray[10][167], dotarray[11][167], dotarray[12][167], dotarray[13][167], dotarray[14][167], dotarray[15][167], dotarray[16][167], dotarray[17][167], dotarray[18][167], dotarray[19][167], dotarray[20][167], dotarray[21][167], dotarray[22][167], dotarray[23][167], dotarray[24][167], dotarray[25][167], dotarray[26][167], dotarray[27][167], dotarray[28][167], dotarray[29][167], dotarray[30][167], dotarray[31][167], dotarray[32][167], dotarray[33][167], dotarray[34][167], dotarray[35][167], dotarray[36][167], dotarray[37][167], dotarray[38][167], dotarray[39][167], dotarray[40][167], dotarray[41][167], dotarray[42][167], dotarray[43][167], dotarray[44][167], dotarray[45][167], dotarray[46][167], dotarray[47][167], dotarray[48][167], dotarray[49][167], dotarray[50][167], dotarray[51][167], dotarray[52][167], dotarray[53][167], dotarray[54][167], dotarray[55][167], dotarray[56][167], dotarray[57][167], dotarray[58][167], dotarray[59][167], dotarray[60][167], dotarray[61][167], dotarray[62][167], dotarray[63][167], dotarray[64][167], dotarray[65][167], dotarray[66][167], dotarray[67][167], dotarray[68][167], dotarray[69][167], dotarray[70][167], dotarray[71][167], dotarray[72][167], dotarray[73][167], dotarray[74][167], dotarray[75][167], dotarray[76][167], dotarray[77][167], dotarray[78][167], dotarray[79][167], dotarray[80][167], dotarray[81][167], dotarray[82][167], dotarray[83][167], dotarray[84][167], dotarray[85][167], dotarray[86][167], dotarray[87][167], dotarray[88][167], dotarray[89][167], dotarray[90][167], dotarray[91][167], dotarray[92][167], dotarray[93][167], dotarray[94][167], dotarray[95][167], dotarray[96][167], dotarray[97][167], dotarray[98][167], dotarray[99][167], dotarray[100][167], dotarray[101][167], dotarray[102][167], dotarray[103][167], dotarray[104][167], dotarray[105][167], dotarray[106][167], dotarray[107][167], dotarray[108][167], dotarray[109][167], dotarray[110][167], dotarray[111][167], dotarray[112][167], dotarray[113][167], dotarray[114][167], dotarray[115][167], dotarray[116][167], dotarray[117][167], dotarray[118][167], dotarray[119][167], dotarray[120][167], dotarray[121][167], dotarray[122][167], dotarray[123][167], dotarray[124][167], dotarray[125][167], dotarray[126][167], dotarray[127][167]};
assign dot_col_168 = {dotarray[0][168], dotarray[1][168], dotarray[2][168], dotarray[3][168], dotarray[4][168], dotarray[5][168], dotarray[6][168], dotarray[7][168], dotarray[8][168], dotarray[9][168], dotarray[10][168], dotarray[11][168], dotarray[12][168], dotarray[13][168], dotarray[14][168], dotarray[15][168], dotarray[16][168], dotarray[17][168], dotarray[18][168], dotarray[19][168], dotarray[20][168], dotarray[21][168], dotarray[22][168], dotarray[23][168], dotarray[24][168], dotarray[25][168], dotarray[26][168], dotarray[27][168], dotarray[28][168], dotarray[29][168], dotarray[30][168], dotarray[31][168], dotarray[32][168], dotarray[33][168], dotarray[34][168], dotarray[35][168], dotarray[36][168], dotarray[37][168], dotarray[38][168], dotarray[39][168], dotarray[40][168], dotarray[41][168], dotarray[42][168], dotarray[43][168], dotarray[44][168], dotarray[45][168], dotarray[46][168], dotarray[47][168], dotarray[48][168], dotarray[49][168], dotarray[50][168], dotarray[51][168], dotarray[52][168], dotarray[53][168], dotarray[54][168], dotarray[55][168], dotarray[56][168], dotarray[57][168], dotarray[58][168], dotarray[59][168], dotarray[60][168], dotarray[61][168], dotarray[62][168], dotarray[63][168], dotarray[64][168], dotarray[65][168], dotarray[66][168], dotarray[67][168], dotarray[68][168], dotarray[69][168], dotarray[70][168], dotarray[71][168], dotarray[72][168], dotarray[73][168], dotarray[74][168], dotarray[75][168], dotarray[76][168], dotarray[77][168], dotarray[78][168], dotarray[79][168], dotarray[80][168], dotarray[81][168], dotarray[82][168], dotarray[83][168], dotarray[84][168], dotarray[85][168], dotarray[86][168], dotarray[87][168], dotarray[88][168], dotarray[89][168], dotarray[90][168], dotarray[91][168], dotarray[92][168], dotarray[93][168], dotarray[94][168], dotarray[95][168], dotarray[96][168], dotarray[97][168], dotarray[98][168], dotarray[99][168], dotarray[100][168], dotarray[101][168], dotarray[102][168], dotarray[103][168], dotarray[104][168], dotarray[105][168], dotarray[106][168], dotarray[107][168], dotarray[108][168], dotarray[109][168], dotarray[110][168], dotarray[111][168], dotarray[112][168], dotarray[113][168], dotarray[114][168], dotarray[115][168], dotarray[116][168], dotarray[117][168], dotarray[118][168], dotarray[119][168], dotarray[120][168], dotarray[121][168], dotarray[122][168], dotarray[123][168], dotarray[124][168], dotarray[125][168], dotarray[126][168], dotarray[127][168]};
assign dot_col_169 = {dotarray[0][169], dotarray[1][169], dotarray[2][169], dotarray[3][169], dotarray[4][169], dotarray[5][169], dotarray[6][169], dotarray[7][169], dotarray[8][169], dotarray[9][169], dotarray[10][169], dotarray[11][169], dotarray[12][169], dotarray[13][169], dotarray[14][169], dotarray[15][169], dotarray[16][169], dotarray[17][169], dotarray[18][169], dotarray[19][169], dotarray[20][169], dotarray[21][169], dotarray[22][169], dotarray[23][169], dotarray[24][169], dotarray[25][169], dotarray[26][169], dotarray[27][169], dotarray[28][169], dotarray[29][169], dotarray[30][169], dotarray[31][169], dotarray[32][169], dotarray[33][169], dotarray[34][169], dotarray[35][169], dotarray[36][169], dotarray[37][169], dotarray[38][169], dotarray[39][169], dotarray[40][169], dotarray[41][169], dotarray[42][169], dotarray[43][169], dotarray[44][169], dotarray[45][169], dotarray[46][169], dotarray[47][169], dotarray[48][169], dotarray[49][169], dotarray[50][169], dotarray[51][169], dotarray[52][169], dotarray[53][169], dotarray[54][169], dotarray[55][169], dotarray[56][169], dotarray[57][169], dotarray[58][169], dotarray[59][169], dotarray[60][169], dotarray[61][169], dotarray[62][169], dotarray[63][169], dotarray[64][169], dotarray[65][169], dotarray[66][169], dotarray[67][169], dotarray[68][169], dotarray[69][169], dotarray[70][169], dotarray[71][169], dotarray[72][169], dotarray[73][169], dotarray[74][169], dotarray[75][169], dotarray[76][169], dotarray[77][169], dotarray[78][169], dotarray[79][169], dotarray[80][169], dotarray[81][169], dotarray[82][169], dotarray[83][169], dotarray[84][169], dotarray[85][169], dotarray[86][169], dotarray[87][169], dotarray[88][169], dotarray[89][169], dotarray[90][169], dotarray[91][169], dotarray[92][169], dotarray[93][169], dotarray[94][169], dotarray[95][169], dotarray[96][169], dotarray[97][169], dotarray[98][169], dotarray[99][169], dotarray[100][169], dotarray[101][169], dotarray[102][169], dotarray[103][169], dotarray[104][169], dotarray[105][169], dotarray[106][169], dotarray[107][169], dotarray[108][169], dotarray[109][169], dotarray[110][169], dotarray[111][169], dotarray[112][169], dotarray[113][169], dotarray[114][169], dotarray[115][169], dotarray[116][169], dotarray[117][169], dotarray[118][169], dotarray[119][169], dotarray[120][169], dotarray[121][169], dotarray[122][169], dotarray[123][169], dotarray[124][169], dotarray[125][169], dotarray[126][169], dotarray[127][169]};
assign dot_col_170 = {dotarray[0][170], dotarray[1][170], dotarray[2][170], dotarray[3][170], dotarray[4][170], dotarray[5][170], dotarray[6][170], dotarray[7][170], dotarray[8][170], dotarray[9][170], dotarray[10][170], dotarray[11][170], dotarray[12][170], dotarray[13][170], dotarray[14][170], dotarray[15][170], dotarray[16][170], dotarray[17][170], dotarray[18][170], dotarray[19][170], dotarray[20][170], dotarray[21][170], dotarray[22][170], dotarray[23][170], dotarray[24][170], dotarray[25][170], dotarray[26][170], dotarray[27][170], dotarray[28][170], dotarray[29][170], dotarray[30][170], dotarray[31][170], dotarray[32][170], dotarray[33][170], dotarray[34][170], dotarray[35][170], dotarray[36][170], dotarray[37][170], dotarray[38][170], dotarray[39][170], dotarray[40][170], dotarray[41][170], dotarray[42][170], dotarray[43][170], dotarray[44][170], dotarray[45][170], dotarray[46][170], dotarray[47][170], dotarray[48][170], dotarray[49][170], dotarray[50][170], dotarray[51][170], dotarray[52][170], dotarray[53][170], dotarray[54][170], dotarray[55][170], dotarray[56][170], dotarray[57][170], dotarray[58][170], dotarray[59][170], dotarray[60][170], dotarray[61][170], dotarray[62][170], dotarray[63][170], dotarray[64][170], dotarray[65][170], dotarray[66][170], dotarray[67][170], dotarray[68][170], dotarray[69][170], dotarray[70][170], dotarray[71][170], dotarray[72][170], dotarray[73][170], dotarray[74][170], dotarray[75][170], dotarray[76][170], dotarray[77][170], dotarray[78][170], dotarray[79][170], dotarray[80][170], dotarray[81][170], dotarray[82][170], dotarray[83][170], dotarray[84][170], dotarray[85][170], dotarray[86][170], dotarray[87][170], dotarray[88][170], dotarray[89][170], dotarray[90][170], dotarray[91][170], dotarray[92][170], dotarray[93][170], dotarray[94][170], dotarray[95][170], dotarray[96][170], dotarray[97][170], dotarray[98][170], dotarray[99][170], dotarray[100][170], dotarray[101][170], dotarray[102][170], dotarray[103][170], dotarray[104][170], dotarray[105][170], dotarray[106][170], dotarray[107][170], dotarray[108][170], dotarray[109][170], dotarray[110][170], dotarray[111][170], dotarray[112][170], dotarray[113][170], dotarray[114][170], dotarray[115][170], dotarray[116][170], dotarray[117][170], dotarray[118][170], dotarray[119][170], dotarray[120][170], dotarray[121][170], dotarray[122][170], dotarray[123][170], dotarray[124][170], dotarray[125][170], dotarray[126][170], dotarray[127][170]};
assign dot_col_171 = {dotarray[0][171], dotarray[1][171], dotarray[2][171], dotarray[3][171], dotarray[4][171], dotarray[5][171], dotarray[6][171], dotarray[7][171], dotarray[8][171], dotarray[9][171], dotarray[10][171], dotarray[11][171], dotarray[12][171], dotarray[13][171], dotarray[14][171], dotarray[15][171], dotarray[16][171], dotarray[17][171], dotarray[18][171], dotarray[19][171], dotarray[20][171], dotarray[21][171], dotarray[22][171], dotarray[23][171], dotarray[24][171], dotarray[25][171], dotarray[26][171], dotarray[27][171], dotarray[28][171], dotarray[29][171], dotarray[30][171], dotarray[31][171], dotarray[32][171], dotarray[33][171], dotarray[34][171], dotarray[35][171], dotarray[36][171], dotarray[37][171], dotarray[38][171], dotarray[39][171], dotarray[40][171], dotarray[41][171], dotarray[42][171], dotarray[43][171], dotarray[44][171], dotarray[45][171], dotarray[46][171], dotarray[47][171], dotarray[48][171], dotarray[49][171], dotarray[50][171], dotarray[51][171], dotarray[52][171], dotarray[53][171], dotarray[54][171], dotarray[55][171], dotarray[56][171], dotarray[57][171], dotarray[58][171], dotarray[59][171], dotarray[60][171], dotarray[61][171], dotarray[62][171], dotarray[63][171], dotarray[64][171], dotarray[65][171], dotarray[66][171], dotarray[67][171], dotarray[68][171], dotarray[69][171], dotarray[70][171], dotarray[71][171], dotarray[72][171], dotarray[73][171], dotarray[74][171], dotarray[75][171], dotarray[76][171], dotarray[77][171], dotarray[78][171], dotarray[79][171], dotarray[80][171], dotarray[81][171], dotarray[82][171], dotarray[83][171], dotarray[84][171], dotarray[85][171], dotarray[86][171], dotarray[87][171], dotarray[88][171], dotarray[89][171], dotarray[90][171], dotarray[91][171], dotarray[92][171], dotarray[93][171], dotarray[94][171], dotarray[95][171], dotarray[96][171], dotarray[97][171], dotarray[98][171], dotarray[99][171], dotarray[100][171], dotarray[101][171], dotarray[102][171], dotarray[103][171], dotarray[104][171], dotarray[105][171], dotarray[106][171], dotarray[107][171], dotarray[108][171], dotarray[109][171], dotarray[110][171], dotarray[111][171], dotarray[112][171], dotarray[113][171], dotarray[114][171], dotarray[115][171], dotarray[116][171], dotarray[117][171], dotarray[118][171], dotarray[119][171], dotarray[120][171], dotarray[121][171], dotarray[122][171], dotarray[123][171], dotarray[124][171], dotarray[125][171], dotarray[126][171], dotarray[127][171]};
assign dot_col_172 = {dotarray[0][172], dotarray[1][172], dotarray[2][172], dotarray[3][172], dotarray[4][172], dotarray[5][172], dotarray[6][172], dotarray[7][172], dotarray[8][172], dotarray[9][172], dotarray[10][172], dotarray[11][172], dotarray[12][172], dotarray[13][172], dotarray[14][172], dotarray[15][172], dotarray[16][172], dotarray[17][172], dotarray[18][172], dotarray[19][172], dotarray[20][172], dotarray[21][172], dotarray[22][172], dotarray[23][172], dotarray[24][172], dotarray[25][172], dotarray[26][172], dotarray[27][172], dotarray[28][172], dotarray[29][172], dotarray[30][172], dotarray[31][172], dotarray[32][172], dotarray[33][172], dotarray[34][172], dotarray[35][172], dotarray[36][172], dotarray[37][172], dotarray[38][172], dotarray[39][172], dotarray[40][172], dotarray[41][172], dotarray[42][172], dotarray[43][172], dotarray[44][172], dotarray[45][172], dotarray[46][172], dotarray[47][172], dotarray[48][172], dotarray[49][172], dotarray[50][172], dotarray[51][172], dotarray[52][172], dotarray[53][172], dotarray[54][172], dotarray[55][172], dotarray[56][172], dotarray[57][172], dotarray[58][172], dotarray[59][172], dotarray[60][172], dotarray[61][172], dotarray[62][172], dotarray[63][172], dotarray[64][172], dotarray[65][172], dotarray[66][172], dotarray[67][172], dotarray[68][172], dotarray[69][172], dotarray[70][172], dotarray[71][172], dotarray[72][172], dotarray[73][172], dotarray[74][172], dotarray[75][172], dotarray[76][172], dotarray[77][172], dotarray[78][172], dotarray[79][172], dotarray[80][172], dotarray[81][172], dotarray[82][172], dotarray[83][172], dotarray[84][172], dotarray[85][172], dotarray[86][172], dotarray[87][172], dotarray[88][172], dotarray[89][172], dotarray[90][172], dotarray[91][172], dotarray[92][172], dotarray[93][172], dotarray[94][172], dotarray[95][172], dotarray[96][172], dotarray[97][172], dotarray[98][172], dotarray[99][172], dotarray[100][172], dotarray[101][172], dotarray[102][172], dotarray[103][172], dotarray[104][172], dotarray[105][172], dotarray[106][172], dotarray[107][172], dotarray[108][172], dotarray[109][172], dotarray[110][172], dotarray[111][172], dotarray[112][172], dotarray[113][172], dotarray[114][172], dotarray[115][172], dotarray[116][172], dotarray[117][172], dotarray[118][172], dotarray[119][172], dotarray[120][172], dotarray[121][172], dotarray[122][172], dotarray[123][172], dotarray[124][172], dotarray[125][172], dotarray[126][172], dotarray[127][172]};
assign dot_col_173 = {dotarray[0][173], dotarray[1][173], dotarray[2][173], dotarray[3][173], dotarray[4][173], dotarray[5][173], dotarray[6][173], dotarray[7][173], dotarray[8][173], dotarray[9][173], dotarray[10][173], dotarray[11][173], dotarray[12][173], dotarray[13][173], dotarray[14][173], dotarray[15][173], dotarray[16][173], dotarray[17][173], dotarray[18][173], dotarray[19][173], dotarray[20][173], dotarray[21][173], dotarray[22][173], dotarray[23][173], dotarray[24][173], dotarray[25][173], dotarray[26][173], dotarray[27][173], dotarray[28][173], dotarray[29][173], dotarray[30][173], dotarray[31][173], dotarray[32][173], dotarray[33][173], dotarray[34][173], dotarray[35][173], dotarray[36][173], dotarray[37][173], dotarray[38][173], dotarray[39][173], dotarray[40][173], dotarray[41][173], dotarray[42][173], dotarray[43][173], dotarray[44][173], dotarray[45][173], dotarray[46][173], dotarray[47][173], dotarray[48][173], dotarray[49][173], dotarray[50][173], dotarray[51][173], dotarray[52][173], dotarray[53][173], dotarray[54][173], dotarray[55][173], dotarray[56][173], dotarray[57][173], dotarray[58][173], dotarray[59][173], dotarray[60][173], dotarray[61][173], dotarray[62][173], dotarray[63][173], dotarray[64][173], dotarray[65][173], dotarray[66][173], dotarray[67][173], dotarray[68][173], dotarray[69][173], dotarray[70][173], dotarray[71][173], dotarray[72][173], dotarray[73][173], dotarray[74][173], dotarray[75][173], dotarray[76][173], dotarray[77][173], dotarray[78][173], dotarray[79][173], dotarray[80][173], dotarray[81][173], dotarray[82][173], dotarray[83][173], dotarray[84][173], dotarray[85][173], dotarray[86][173], dotarray[87][173], dotarray[88][173], dotarray[89][173], dotarray[90][173], dotarray[91][173], dotarray[92][173], dotarray[93][173], dotarray[94][173], dotarray[95][173], dotarray[96][173], dotarray[97][173], dotarray[98][173], dotarray[99][173], dotarray[100][173], dotarray[101][173], dotarray[102][173], dotarray[103][173], dotarray[104][173], dotarray[105][173], dotarray[106][173], dotarray[107][173], dotarray[108][173], dotarray[109][173], dotarray[110][173], dotarray[111][173], dotarray[112][173], dotarray[113][173], dotarray[114][173], dotarray[115][173], dotarray[116][173], dotarray[117][173], dotarray[118][173], dotarray[119][173], dotarray[120][173], dotarray[121][173], dotarray[122][173], dotarray[123][173], dotarray[124][173], dotarray[125][173], dotarray[126][173], dotarray[127][173]};
assign dot_col_174 = {dotarray[0][174], dotarray[1][174], dotarray[2][174], dotarray[3][174], dotarray[4][174], dotarray[5][174], dotarray[6][174], dotarray[7][174], dotarray[8][174], dotarray[9][174], dotarray[10][174], dotarray[11][174], dotarray[12][174], dotarray[13][174], dotarray[14][174], dotarray[15][174], dotarray[16][174], dotarray[17][174], dotarray[18][174], dotarray[19][174], dotarray[20][174], dotarray[21][174], dotarray[22][174], dotarray[23][174], dotarray[24][174], dotarray[25][174], dotarray[26][174], dotarray[27][174], dotarray[28][174], dotarray[29][174], dotarray[30][174], dotarray[31][174], dotarray[32][174], dotarray[33][174], dotarray[34][174], dotarray[35][174], dotarray[36][174], dotarray[37][174], dotarray[38][174], dotarray[39][174], dotarray[40][174], dotarray[41][174], dotarray[42][174], dotarray[43][174], dotarray[44][174], dotarray[45][174], dotarray[46][174], dotarray[47][174], dotarray[48][174], dotarray[49][174], dotarray[50][174], dotarray[51][174], dotarray[52][174], dotarray[53][174], dotarray[54][174], dotarray[55][174], dotarray[56][174], dotarray[57][174], dotarray[58][174], dotarray[59][174], dotarray[60][174], dotarray[61][174], dotarray[62][174], dotarray[63][174], dotarray[64][174], dotarray[65][174], dotarray[66][174], dotarray[67][174], dotarray[68][174], dotarray[69][174], dotarray[70][174], dotarray[71][174], dotarray[72][174], dotarray[73][174], dotarray[74][174], dotarray[75][174], dotarray[76][174], dotarray[77][174], dotarray[78][174], dotarray[79][174], dotarray[80][174], dotarray[81][174], dotarray[82][174], dotarray[83][174], dotarray[84][174], dotarray[85][174], dotarray[86][174], dotarray[87][174], dotarray[88][174], dotarray[89][174], dotarray[90][174], dotarray[91][174], dotarray[92][174], dotarray[93][174], dotarray[94][174], dotarray[95][174], dotarray[96][174], dotarray[97][174], dotarray[98][174], dotarray[99][174], dotarray[100][174], dotarray[101][174], dotarray[102][174], dotarray[103][174], dotarray[104][174], dotarray[105][174], dotarray[106][174], dotarray[107][174], dotarray[108][174], dotarray[109][174], dotarray[110][174], dotarray[111][174], dotarray[112][174], dotarray[113][174], dotarray[114][174], dotarray[115][174], dotarray[116][174], dotarray[117][174], dotarray[118][174], dotarray[119][174], dotarray[120][174], dotarray[121][174], dotarray[122][174], dotarray[123][174], dotarray[124][174], dotarray[125][174], dotarray[126][174], dotarray[127][174]};
assign dot_col_175 = {dotarray[0][175], dotarray[1][175], dotarray[2][175], dotarray[3][175], dotarray[4][175], dotarray[5][175], dotarray[6][175], dotarray[7][175], dotarray[8][175], dotarray[9][175], dotarray[10][175], dotarray[11][175], dotarray[12][175], dotarray[13][175], dotarray[14][175], dotarray[15][175], dotarray[16][175], dotarray[17][175], dotarray[18][175], dotarray[19][175], dotarray[20][175], dotarray[21][175], dotarray[22][175], dotarray[23][175], dotarray[24][175], dotarray[25][175], dotarray[26][175], dotarray[27][175], dotarray[28][175], dotarray[29][175], dotarray[30][175], dotarray[31][175], dotarray[32][175], dotarray[33][175], dotarray[34][175], dotarray[35][175], dotarray[36][175], dotarray[37][175], dotarray[38][175], dotarray[39][175], dotarray[40][175], dotarray[41][175], dotarray[42][175], dotarray[43][175], dotarray[44][175], dotarray[45][175], dotarray[46][175], dotarray[47][175], dotarray[48][175], dotarray[49][175], dotarray[50][175], dotarray[51][175], dotarray[52][175], dotarray[53][175], dotarray[54][175], dotarray[55][175], dotarray[56][175], dotarray[57][175], dotarray[58][175], dotarray[59][175], dotarray[60][175], dotarray[61][175], dotarray[62][175], dotarray[63][175], dotarray[64][175], dotarray[65][175], dotarray[66][175], dotarray[67][175], dotarray[68][175], dotarray[69][175], dotarray[70][175], dotarray[71][175], dotarray[72][175], dotarray[73][175], dotarray[74][175], dotarray[75][175], dotarray[76][175], dotarray[77][175], dotarray[78][175], dotarray[79][175], dotarray[80][175], dotarray[81][175], dotarray[82][175], dotarray[83][175], dotarray[84][175], dotarray[85][175], dotarray[86][175], dotarray[87][175], dotarray[88][175], dotarray[89][175], dotarray[90][175], dotarray[91][175], dotarray[92][175], dotarray[93][175], dotarray[94][175], dotarray[95][175], dotarray[96][175], dotarray[97][175], dotarray[98][175], dotarray[99][175], dotarray[100][175], dotarray[101][175], dotarray[102][175], dotarray[103][175], dotarray[104][175], dotarray[105][175], dotarray[106][175], dotarray[107][175], dotarray[108][175], dotarray[109][175], dotarray[110][175], dotarray[111][175], dotarray[112][175], dotarray[113][175], dotarray[114][175], dotarray[115][175], dotarray[116][175], dotarray[117][175], dotarray[118][175], dotarray[119][175], dotarray[120][175], dotarray[121][175], dotarray[122][175], dotarray[123][175], dotarray[124][175], dotarray[125][175], dotarray[126][175], dotarray[127][175]};
assign dot_col_176 = {dotarray[0][176], dotarray[1][176], dotarray[2][176], dotarray[3][176], dotarray[4][176], dotarray[5][176], dotarray[6][176], dotarray[7][176], dotarray[8][176], dotarray[9][176], dotarray[10][176], dotarray[11][176], dotarray[12][176], dotarray[13][176], dotarray[14][176], dotarray[15][176], dotarray[16][176], dotarray[17][176], dotarray[18][176], dotarray[19][176], dotarray[20][176], dotarray[21][176], dotarray[22][176], dotarray[23][176], dotarray[24][176], dotarray[25][176], dotarray[26][176], dotarray[27][176], dotarray[28][176], dotarray[29][176], dotarray[30][176], dotarray[31][176], dotarray[32][176], dotarray[33][176], dotarray[34][176], dotarray[35][176], dotarray[36][176], dotarray[37][176], dotarray[38][176], dotarray[39][176], dotarray[40][176], dotarray[41][176], dotarray[42][176], dotarray[43][176], dotarray[44][176], dotarray[45][176], dotarray[46][176], dotarray[47][176], dotarray[48][176], dotarray[49][176], dotarray[50][176], dotarray[51][176], dotarray[52][176], dotarray[53][176], dotarray[54][176], dotarray[55][176], dotarray[56][176], dotarray[57][176], dotarray[58][176], dotarray[59][176], dotarray[60][176], dotarray[61][176], dotarray[62][176], dotarray[63][176], dotarray[64][176], dotarray[65][176], dotarray[66][176], dotarray[67][176], dotarray[68][176], dotarray[69][176], dotarray[70][176], dotarray[71][176], dotarray[72][176], dotarray[73][176], dotarray[74][176], dotarray[75][176], dotarray[76][176], dotarray[77][176], dotarray[78][176], dotarray[79][176], dotarray[80][176], dotarray[81][176], dotarray[82][176], dotarray[83][176], dotarray[84][176], dotarray[85][176], dotarray[86][176], dotarray[87][176], dotarray[88][176], dotarray[89][176], dotarray[90][176], dotarray[91][176], dotarray[92][176], dotarray[93][176], dotarray[94][176], dotarray[95][176], dotarray[96][176], dotarray[97][176], dotarray[98][176], dotarray[99][176], dotarray[100][176], dotarray[101][176], dotarray[102][176], dotarray[103][176], dotarray[104][176], dotarray[105][176], dotarray[106][176], dotarray[107][176], dotarray[108][176], dotarray[109][176], dotarray[110][176], dotarray[111][176], dotarray[112][176], dotarray[113][176], dotarray[114][176], dotarray[115][176], dotarray[116][176], dotarray[117][176], dotarray[118][176], dotarray[119][176], dotarray[120][176], dotarray[121][176], dotarray[122][176], dotarray[123][176], dotarray[124][176], dotarray[125][176], dotarray[126][176], dotarray[127][176]};
assign dot_col_177 = {dotarray[0][177], dotarray[1][177], dotarray[2][177], dotarray[3][177], dotarray[4][177], dotarray[5][177], dotarray[6][177], dotarray[7][177], dotarray[8][177], dotarray[9][177], dotarray[10][177], dotarray[11][177], dotarray[12][177], dotarray[13][177], dotarray[14][177], dotarray[15][177], dotarray[16][177], dotarray[17][177], dotarray[18][177], dotarray[19][177], dotarray[20][177], dotarray[21][177], dotarray[22][177], dotarray[23][177], dotarray[24][177], dotarray[25][177], dotarray[26][177], dotarray[27][177], dotarray[28][177], dotarray[29][177], dotarray[30][177], dotarray[31][177], dotarray[32][177], dotarray[33][177], dotarray[34][177], dotarray[35][177], dotarray[36][177], dotarray[37][177], dotarray[38][177], dotarray[39][177], dotarray[40][177], dotarray[41][177], dotarray[42][177], dotarray[43][177], dotarray[44][177], dotarray[45][177], dotarray[46][177], dotarray[47][177], dotarray[48][177], dotarray[49][177], dotarray[50][177], dotarray[51][177], dotarray[52][177], dotarray[53][177], dotarray[54][177], dotarray[55][177], dotarray[56][177], dotarray[57][177], dotarray[58][177], dotarray[59][177], dotarray[60][177], dotarray[61][177], dotarray[62][177], dotarray[63][177], dotarray[64][177], dotarray[65][177], dotarray[66][177], dotarray[67][177], dotarray[68][177], dotarray[69][177], dotarray[70][177], dotarray[71][177], dotarray[72][177], dotarray[73][177], dotarray[74][177], dotarray[75][177], dotarray[76][177], dotarray[77][177], dotarray[78][177], dotarray[79][177], dotarray[80][177], dotarray[81][177], dotarray[82][177], dotarray[83][177], dotarray[84][177], dotarray[85][177], dotarray[86][177], dotarray[87][177], dotarray[88][177], dotarray[89][177], dotarray[90][177], dotarray[91][177], dotarray[92][177], dotarray[93][177], dotarray[94][177], dotarray[95][177], dotarray[96][177], dotarray[97][177], dotarray[98][177], dotarray[99][177], dotarray[100][177], dotarray[101][177], dotarray[102][177], dotarray[103][177], dotarray[104][177], dotarray[105][177], dotarray[106][177], dotarray[107][177], dotarray[108][177], dotarray[109][177], dotarray[110][177], dotarray[111][177], dotarray[112][177], dotarray[113][177], dotarray[114][177], dotarray[115][177], dotarray[116][177], dotarray[117][177], dotarray[118][177], dotarray[119][177], dotarray[120][177], dotarray[121][177], dotarray[122][177], dotarray[123][177], dotarray[124][177], dotarray[125][177], dotarray[126][177], dotarray[127][177]};
assign dot_col_178 = {dotarray[0][178], dotarray[1][178], dotarray[2][178], dotarray[3][178], dotarray[4][178], dotarray[5][178], dotarray[6][178], dotarray[7][178], dotarray[8][178], dotarray[9][178], dotarray[10][178], dotarray[11][178], dotarray[12][178], dotarray[13][178], dotarray[14][178], dotarray[15][178], dotarray[16][178], dotarray[17][178], dotarray[18][178], dotarray[19][178], dotarray[20][178], dotarray[21][178], dotarray[22][178], dotarray[23][178], dotarray[24][178], dotarray[25][178], dotarray[26][178], dotarray[27][178], dotarray[28][178], dotarray[29][178], dotarray[30][178], dotarray[31][178], dotarray[32][178], dotarray[33][178], dotarray[34][178], dotarray[35][178], dotarray[36][178], dotarray[37][178], dotarray[38][178], dotarray[39][178], dotarray[40][178], dotarray[41][178], dotarray[42][178], dotarray[43][178], dotarray[44][178], dotarray[45][178], dotarray[46][178], dotarray[47][178], dotarray[48][178], dotarray[49][178], dotarray[50][178], dotarray[51][178], dotarray[52][178], dotarray[53][178], dotarray[54][178], dotarray[55][178], dotarray[56][178], dotarray[57][178], dotarray[58][178], dotarray[59][178], dotarray[60][178], dotarray[61][178], dotarray[62][178], dotarray[63][178], dotarray[64][178], dotarray[65][178], dotarray[66][178], dotarray[67][178], dotarray[68][178], dotarray[69][178], dotarray[70][178], dotarray[71][178], dotarray[72][178], dotarray[73][178], dotarray[74][178], dotarray[75][178], dotarray[76][178], dotarray[77][178], dotarray[78][178], dotarray[79][178], dotarray[80][178], dotarray[81][178], dotarray[82][178], dotarray[83][178], dotarray[84][178], dotarray[85][178], dotarray[86][178], dotarray[87][178], dotarray[88][178], dotarray[89][178], dotarray[90][178], dotarray[91][178], dotarray[92][178], dotarray[93][178], dotarray[94][178], dotarray[95][178], dotarray[96][178], dotarray[97][178], dotarray[98][178], dotarray[99][178], dotarray[100][178], dotarray[101][178], dotarray[102][178], dotarray[103][178], dotarray[104][178], dotarray[105][178], dotarray[106][178], dotarray[107][178], dotarray[108][178], dotarray[109][178], dotarray[110][178], dotarray[111][178], dotarray[112][178], dotarray[113][178], dotarray[114][178], dotarray[115][178], dotarray[116][178], dotarray[117][178], dotarray[118][178], dotarray[119][178], dotarray[120][178], dotarray[121][178], dotarray[122][178], dotarray[123][178], dotarray[124][178], dotarray[125][178], dotarray[126][178], dotarray[127][178]};
assign dot_col_179 = {dotarray[0][179], dotarray[1][179], dotarray[2][179], dotarray[3][179], dotarray[4][179], dotarray[5][179], dotarray[6][179], dotarray[7][179], dotarray[8][179], dotarray[9][179], dotarray[10][179], dotarray[11][179], dotarray[12][179], dotarray[13][179], dotarray[14][179], dotarray[15][179], dotarray[16][179], dotarray[17][179], dotarray[18][179], dotarray[19][179], dotarray[20][179], dotarray[21][179], dotarray[22][179], dotarray[23][179], dotarray[24][179], dotarray[25][179], dotarray[26][179], dotarray[27][179], dotarray[28][179], dotarray[29][179], dotarray[30][179], dotarray[31][179], dotarray[32][179], dotarray[33][179], dotarray[34][179], dotarray[35][179], dotarray[36][179], dotarray[37][179], dotarray[38][179], dotarray[39][179], dotarray[40][179], dotarray[41][179], dotarray[42][179], dotarray[43][179], dotarray[44][179], dotarray[45][179], dotarray[46][179], dotarray[47][179], dotarray[48][179], dotarray[49][179], dotarray[50][179], dotarray[51][179], dotarray[52][179], dotarray[53][179], dotarray[54][179], dotarray[55][179], dotarray[56][179], dotarray[57][179], dotarray[58][179], dotarray[59][179], dotarray[60][179], dotarray[61][179], dotarray[62][179], dotarray[63][179], dotarray[64][179], dotarray[65][179], dotarray[66][179], dotarray[67][179], dotarray[68][179], dotarray[69][179], dotarray[70][179], dotarray[71][179], dotarray[72][179], dotarray[73][179], dotarray[74][179], dotarray[75][179], dotarray[76][179], dotarray[77][179], dotarray[78][179], dotarray[79][179], dotarray[80][179], dotarray[81][179], dotarray[82][179], dotarray[83][179], dotarray[84][179], dotarray[85][179], dotarray[86][179], dotarray[87][179], dotarray[88][179], dotarray[89][179], dotarray[90][179], dotarray[91][179], dotarray[92][179], dotarray[93][179], dotarray[94][179], dotarray[95][179], dotarray[96][179], dotarray[97][179], dotarray[98][179], dotarray[99][179], dotarray[100][179], dotarray[101][179], dotarray[102][179], dotarray[103][179], dotarray[104][179], dotarray[105][179], dotarray[106][179], dotarray[107][179], dotarray[108][179], dotarray[109][179], dotarray[110][179], dotarray[111][179], dotarray[112][179], dotarray[113][179], dotarray[114][179], dotarray[115][179], dotarray[116][179], dotarray[117][179], dotarray[118][179], dotarray[119][179], dotarray[120][179], dotarray[121][179], dotarray[122][179], dotarray[123][179], dotarray[124][179], dotarray[125][179], dotarray[126][179], dotarray[127][179]};
assign dot_col_180 = {dotarray[0][180], dotarray[1][180], dotarray[2][180], dotarray[3][180], dotarray[4][180], dotarray[5][180], dotarray[6][180], dotarray[7][180], dotarray[8][180], dotarray[9][180], dotarray[10][180], dotarray[11][180], dotarray[12][180], dotarray[13][180], dotarray[14][180], dotarray[15][180], dotarray[16][180], dotarray[17][180], dotarray[18][180], dotarray[19][180], dotarray[20][180], dotarray[21][180], dotarray[22][180], dotarray[23][180], dotarray[24][180], dotarray[25][180], dotarray[26][180], dotarray[27][180], dotarray[28][180], dotarray[29][180], dotarray[30][180], dotarray[31][180], dotarray[32][180], dotarray[33][180], dotarray[34][180], dotarray[35][180], dotarray[36][180], dotarray[37][180], dotarray[38][180], dotarray[39][180], dotarray[40][180], dotarray[41][180], dotarray[42][180], dotarray[43][180], dotarray[44][180], dotarray[45][180], dotarray[46][180], dotarray[47][180], dotarray[48][180], dotarray[49][180], dotarray[50][180], dotarray[51][180], dotarray[52][180], dotarray[53][180], dotarray[54][180], dotarray[55][180], dotarray[56][180], dotarray[57][180], dotarray[58][180], dotarray[59][180], dotarray[60][180], dotarray[61][180], dotarray[62][180], dotarray[63][180], dotarray[64][180], dotarray[65][180], dotarray[66][180], dotarray[67][180], dotarray[68][180], dotarray[69][180], dotarray[70][180], dotarray[71][180], dotarray[72][180], dotarray[73][180], dotarray[74][180], dotarray[75][180], dotarray[76][180], dotarray[77][180], dotarray[78][180], dotarray[79][180], dotarray[80][180], dotarray[81][180], dotarray[82][180], dotarray[83][180], dotarray[84][180], dotarray[85][180], dotarray[86][180], dotarray[87][180], dotarray[88][180], dotarray[89][180], dotarray[90][180], dotarray[91][180], dotarray[92][180], dotarray[93][180], dotarray[94][180], dotarray[95][180], dotarray[96][180], dotarray[97][180], dotarray[98][180], dotarray[99][180], dotarray[100][180], dotarray[101][180], dotarray[102][180], dotarray[103][180], dotarray[104][180], dotarray[105][180], dotarray[106][180], dotarray[107][180], dotarray[108][180], dotarray[109][180], dotarray[110][180], dotarray[111][180], dotarray[112][180], dotarray[113][180], dotarray[114][180], dotarray[115][180], dotarray[116][180], dotarray[117][180], dotarray[118][180], dotarray[119][180], dotarray[120][180], dotarray[121][180], dotarray[122][180], dotarray[123][180], dotarray[124][180], dotarray[125][180], dotarray[126][180], dotarray[127][180]};
assign dot_col_181 = {dotarray[0][181], dotarray[1][181], dotarray[2][181], dotarray[3][181], dotarray[4][181], dotarray[5][181], dotarray[6][181], dotarray[7][181], dotarray[8][181], dotarray[9][181], dotarray[10][181], dotarray[11][181], dotarray[12][181], dotarray[13][181], dotarray[14][181], dotarray[15][181], dotarray[16][181], dotarray[17][181], dotarray[18][181], dotarray[19][181], dotarray[20][181], dotarray[21][181], dotarray[22][181], dotarray[23][181], dotarray[24][181], dotarray[25][181], dotarray[26][181], dotarray[27][181], dotarray[28][181], dotarray[29][181], dotarray[30][181], dotarray[31][181], dotarray[32][181], dotarray[33][181], dotarray[34][181], dotarray[35][181], dotarray[36][181], dotarray[37][181], dotarray[38][181], dotarray[39][181], dotarray[40][181], dotarray[41][181], dotarray[42][181], dotarray[43][181], dotarray[44][181], dotarray[45][181], dotarray[46][181], dotarray[47][181], dotarray[48][181], dotarray[49][181], dotarray[50][181], dotarray[51][181], dotarray[52][181], dotarray[53][181], dotarray[54][181], dotarray[55][181], dotarray[56][181], dotarray[57][181], dotarray[58][181], dotarray[59][181], dotarray[60][181], dotarray[61][181], dotarray[62][181], dotarray[63][181], dotarray[64][181], dotarray[65][181], dotarray[66][181], dotarray[67][181], dotarray[68][181], dotarray[69][181], dotarray[70][181], dotarray[71][181], dotarray[72][181], dotarray[73][181], dotarray[74][181], dotarray[75][181], dotarray[76][181], dotarray[77][181], dotarray[78][181], dotarray[79][181], dotarray[80][181], dotarray[81][181], dotarray[82][181], dotarray[83][181], dotarray[84][181], dotarray[85][181], dotarray[86][181], dotarray[87][181], dotarray[88][181], dotarray[89][181], dotarray[90][181], dotarray[91][181], dotarray[92][181], dotarray[93][181], dotarray[94][181], dotarray[95][181], dotarray[96][181], dotarray[97][181], dotarray[98][181], dotarray[99][181], dotarray[100][181], dotarray[101][181], dotarray[102][181], dotarray[103][181], dotarray[104][181], dotarray[105][181], dotarray[106][181], dotarray[107][181], dotarray[108][181], dotarray[109][181], dotarray[110][181], dotarray[111][181], dotarray[112][181], dotarray[113][181], dotarray[114][181], dotarray[115][181], dotarray[116][181], dotarray[117][181], dotarray[118][181], dotarray[119][181], dotarray[120][181], dotarray[121][181], dotarray[122][181], dotarray[123][181], dotarray[124][181], dotarray[125][181], dotarray[126][181], dotarray[127][181]};
assign dot_col_182 = {dotarray[0][182], dotarray[1][182], dotarray[2][182], dotarray[3][182], dotarray[4][182], dotarray[5][182], dotarray[6][182], dotarray[7][182], dotarray[8][182], dotarray[9][182], dotarray[10][182], dotarray[11][182], dotarray[12][182], dotarray[13][182], dotarray[14][182], dotarray[15][182], dotarray[16][182], dotarray[17][182], dotarray[18][182], dotarray[19][182], dotarray[20][182], dotarray[21][182], dotarray[22][182], dotarray[23][182], dotarray[24][182], dotarray[25][182], dotarray[26][182], dotarray[27][182], dotarray[28][182], dotarray[29][182], dotarray[30][182], dotarray[31][182], dotarray[32][182], dotarray[33][182], dotarray[34][182], dotarray[35][182], dotarray[36][182], dotarray[37][182], dotarray[38][182], dotarray[39][182], dotarray[40][182], dotarray[41][182], dotarray[42][182], dotarray[43][182], dotarray[44][182], dotarray[45][182], dotarray[46][182], dotarray[47][182], dotarray[48][182], dotarray[49][182], dotarray[50][182], dotarray[51][182], dotarray[52][182], dotarray[53][182], dotarray[54][182], dotarray[55][182], dotarray[56][182], dotarray[57][182], dotarray[58][182], dotarray[59][182], dotarray[60][182], dotarray[61][182], dotarray[62][182], dotarray[63][182], dotarray[64][182], dotarray[65][182], dotarray[66][182], dotarray[67][182], dotarray[68][182], dotarray[69][182], dotarray[70][182], dotarray[71][182], dotarray[72][182], dotarray[73][182], dotarray[74][182], dotarray[75][182], dotarray[76][182], dotarray[77][182], dotarray[78][182], dotarray[79][182], dotarray[80][182], dotarray[81][182], dotarray[82][182], dotarray[83][182], dotarray[84][182], dotarray[85][182], dotarray[86][182], dotarray[87][182], dotarray[88][182], dotarray[89][182], dotarray[90][182], dotarray[91][182], dotarray[92][182], dotarray[93][182], dotarray[94][182], dotarray[95][182], dotarray[96][182], dotarray[97][182], dotarray[98][182], dotarray[99][182], dotarray[100][182], dotarray[101][182], dotarray[102][182], dotarray[103][182], dotarray[104][182], dotarray[105][182], dotarray[106][182], dotarray[107][182], dotarray[108][182], dotarray[109][182], dotarray[110][182], dotarray[111][182], dotarray[112][182], dotarray[113][182], dotarray[114][182], dotarray[115][182], dotarray[116][182], dotarray[117][182], dotarray[118][182], dotarray[119][182], dotarray[120][182], dotarray[121][182], dotarray[122][182], dotarray[123][182], dotarray[124][182], dotarray[125][182], dotarray[126][182], dotarray[127][182]};
assign dot_col_183 = {dotarray[0][183], dotarray[1][183], dotarray[2][183], dotarray[3][183], dotarray[4][183], dotarray[5][183], dotarray[6][183], dotarray[7][183], dotarray[8][183], dotarray[9][183], dotarray[10][183], dotarray[11][183], dotarray[12][183], dotarray[13][183], dotarray[14][183], dotarray[15][183], dotarray[16][183], dotarray[17][183], dotarray[18][183], dotarray[19][183], dotarray[20][183], dotarray[21][183], dotarray[22][183], dotarray[23][183], dotarray[24][183], dotarray[25][183], dotarray[26][183], dotarray[27][183], dotarray[28][183], dotarray[29][183], dotarray[30][183], dotarray[31][183], dotarray[32][183], dotarray[33][183], dotarray[34][183], dotarray[35][183], dotarray[36][183], dotarray[37][183], dotarray[38][183], dotarray[39][183], dotarray[40][183], dotarray[41][183], dotarray[42][183], dotarray[43][183], dotarray[44][183], dotarray[45][183], dotarray[46][183], dotarray[47][183], dotarray[48][183], dotarray[49][183], dotarray[50][183], dotarray[51][183], dotarray[52][183], dotarray[53][183], dotarray[54][183], dotarray[55][183], dotarray[56][183], dotarray[57][183], dotarray[58][183], dotarray[59][183], dotarray[60][183], dotarray[61][183], dotarray[62][183], dotarray[63][183], dotarray[64][183], dotarray[65][183], dotarray[66][183], dotarray[67][183], dotarray[68][183], dotarray[69][183], dotarray[70][183], dotarray[71][183], dotarray[72][183], dotarray[73][183], dotarray[74][183], dotarray[75][183], dotarray[76][183], dotarray[77][183], dotarray[78][183], dotarray[79][183], dotarray[80][183], dotarray[81][183], dotarray[82][183], dotarray[83][183], dotarray[84][183], dotarray[85][183], dotarray[86][183], dotarray[87][183], dotarray[88][183], dotarray[89][183], dotarray[90][183], dotarray[91][183], dotarray[92][183], dotarray[93][183], dotarray[94][183], dotarray[95][183], dotarray[96][183], dotarray[97][183], dotarray[98][183], dotarray[99][183], dotarray[100][183], dotarray[101][183], dotarray[102][183], dotarray[103][183], dotarray[104][183], dotarray[105][183], dotarray[106][183], dotarray[107][183], dotarray[108][183], dotarray[109][183], dotarray[110][183], dotarray[111][183], dotarray[112][183], dotarray[113][183], dotarray[114][183], dotarray[115][183], dotarray[116][183], dotarray[117][183], dotarray[118][183], dotarray[119][183], dotarray[120][183], dotarray[121][183], dotarray[122][183], dotarray[123][183], dotarray[124][183], dotarray[125][183], dotarray[126][183], dotarray[127][183]};
assign dot_col_184 = {dotarray[0][184], dotarray[1][184], dotarray[2][184], dotarray[3][184], dotarray[4][184], dotarray[5][184], dotarray[6][184], dotarray[7][184], dotarray[8][184], dotarray[9][184], dotarray[10][184], dotarray[11][184], dotarray[12][184], dotarray[13][184], dotarray[14][184], dotarray[15][184], dotarray[16][184], dotarray[17][184], dotarray[18][184], dotarray[19][184], dotarray[20][184], dotarray[21][184], dotarray[22][184], dotarray[23][184], dotarray[24][184], dotarray[25][184], dotarray[26][184], dotarray[27][184], dotarray[28][184], dotarray[29][184], dotarray[30][184], dotarray[31][184], dotarray[32][184], dotarray[33][184], dotarray[34][184], dotarray[35][184], dotarray[36][184], dotarray[37][184], dotarray[38][184], dotarray[39][184], dotarray[40][184], dotarray[41][184], dotarray[42][184], dotarray[43][184], dotarray[44][184], dotarray[45][184], dotarray[46][184], dotarray[47][184], dotarray[48][184], dotarray[49][184], dotarray[50][184], dotarray[51][184], dotarray[52][184], dotarray[53][184], dotarray[54][184], dotarray[55][184], dotarray[56][184], dotarray[57][184], dotarray[58][184], dotarray[59][184], dotarray[60][184], dotarray[61][184], dotarray[62][184], dotarray[63][184], dotarray[64][184], dotarray[65][184], dotarray[66][184], dotarray[67][184], dotarray[68][184], dotarray[69][184], dotarray[70][184], dotarray[71][184], dotarray[72][184], dotarray[73][184], dotarray[74][184], dotarray[75][184], dotarray[76][184], dotarray[77][184], dotarray[78][184], dotarray[79][184], dotarray[80][184], dotarray[81][184], dotarray[82][184], dotarray[83][184], dotarray[84][184], dotarray[85][184], dotarray[86][184], dotarray[87][184], dotarray[88][184], dotarray[89][184], dotarray[90][184], dotarray[91][184], dotarray[92][184], dotarray[93][184], dotarray[94][184], dotarray[95][184], dotarray[96][184], dotarray[97][184], dotarray[98][184], dotarray[99][184], dotarray[100][184], dotarray[101][184], dotarray[102][184], dotarray[103][184], dotarray[104][184], dotarray[105][184], dotarray[106][184], dotarray[107][184], dotarray[108][184], dotarray[109][184], dotarray[110][184], dotarray[111][184], dotarray[112][184], dotarray[113][184], dotarray[114][184], dotarray[115][184], dotarray[116][184], dotarray[117][184], dotarray[118][184], dotarray[119][184], dotarray[120][184], dotarray[121][184], dotarray[122][184], dotarray[123][184], dotarray[124][184], dotarray[125][184], dotarray[126][184], dotarray[127][184]};
assign dot_col_185 = {dotarray[0][185], dotarray[1][185], dotarray[2][185], dotarray[3][185], dotarray[4][185], dotarray[5][185], dotarray[6][185], dotarray[7][185], dotarray[8][185], dotarray[9][185], dotarray[10][185], dotarray[11][185], dotarray[12][185], dotarray[13][185], dotarray[14][185], dotarray[15][185], dotarray[16][185], dotarray[17][185], dotarray[18][185], dotarray[19][185], dotarray[20][185], dotarray[21][185], dotarray[22][185], dotarray[23][185], dotarray[24][185], dotarray[25][185], dotarray[26][185], dotarray[27][185], dotarray[28][185], dotarray[29][185], dotarray[30][185], dotarray[31][185], dotarray[32][185], dotarray[33][185], dotarray[34][185], dotarray[35][185], dotarray[36][185], dotarray[37][185], dotarray[38][185], dotarray[39][185], dotarray[40][185], dotarray[41][185], dotarray[42][185], dotarray[43][185], dotarray[44][185], dotarray[45][185], dotarray[46][185], dotarray[47][185], dotarray[48][185], dotarray[49][185], dotarray[50][185], dotarray[51][185], dotarray[52][185], dotarray[53][185], dotarray[54][185], dotarray[55][185], dotarray[56][185], dotarray[57][185], dotarray[58][185], dotarray[59][185], dotarray[60][185], dotarray[61][185], dotarray[62][185], dotarray[63][185], dotarray[64][185], dotarray[65][185], dotarray[66][185], dotarray[67][185], dotarray[68][185], dotarray[69][185], dotarray[70][185], dotarray[71][185], dotarray[72][185], dotarray[73][185], dotarray[74][185], dotarray[75][185], dotarray[76][185], dotarray[77][185], dotarray[78][185], dotarray[79][185], dotarray[80][185], dotarray[81][185], dotarray[82][185], dotarray[83][185], dotarray[84][185], dotarray[85][185], dotarray[86][185], dotarray[87][185], dotarray[88][185], dotarray[89][185], dotarray[90][185], dotarray[91][185], dotarray[92][185], dotarray[93][185], dotarray[94][185], dotarray[95][185], dotarray[96][185], dotarray[97][185], dotarray[98][185], dotarray[99][185], dotarray[100][185], dotarray[101][185], dotarray[102][185], dotarray[103][185], dotarray[104][185], dotarray[105][185], dotarray[106][185], dotarray[107][185], dotarray[108][185], dotarray[109][185], dotarray[110][185], dotarray[111][185], dotarray[112][185], dotarray[113][185], dotarray[114][185], dotarray[115][185], dotarray[116][185], dotarray[117][185], dotarray[118][185], dotarray[119][185], dotarray[120][185], dotarray[121][185], dotarray[122][185], dotarray[123][185], dotarray[124][185], dotarray[125][185], dotarray[126][185], dotarray[127][185]};
assign dot_col_186 = {dotarray[0][186], dotarray[1][186], dotarray[2][186], dotarray[3][186], dotarray[4][186], dotarray[5][186], dotarray[6][186], dotarray[7][186], dotarray[8][186], dotarray[9][186], dotarray[10][186], dotarray[11][186], dotarray[12][186], dotarray[13][186], dotarray[14][186], dotarray[15][186], dotarray[16][186], dotarray[17][186], dotarray[18][186], dotarray[19][186], dotarray[20][186], dotarray[21][186], dotarray[22][186], dotarray[23][186], dotarray[24][186], dotarray[25][186], dotarray[26][186], dotarray[27][186], dotarray[28][186], dotarray[29][186], dotarray[30][186], dotarray[31][186], dotarray[32][186], dotarray[33][186], dotarray[34][186], dotarray[35][186], dotarray[36][186], dotarray[37][186], dotarray[38][186], dotarray[39][186], dotarray[40][186], dotarray[41][186], dotarray[42][186], dotarray[43][186], dotarray[44][186], dotarray[45][186], dotarray[46][186], dotarray[47][186], dotarray[48][186], dotarray[49][186], dotarray[50][186], dotarray[51][186], dotarray[52][186], dotarray[53][186], dotarray[54][186], dotarray[55][186], dotarray[56][186], dotarray[57][186], dotarray[58][186], dotarray[59][186], dotarray[60][186], dotarray[61][186], dotarray[62][186], dotarray[63][186], dotarray[64][186], dotarray[65][186], dotarray[66][186], dotarray[67][186], dotarray[68][186], dotarray[69][186], dotarray[70][186], dotarray[71][186], dotarray[72][186], dotarray[73][186], dotarray[74][186], dotarray[75][186], dotarray[76][186], dotarray[77][186], dotarray[78][186], dotarray[79][186], dotarray[80][186], dotarray[81][186], dotarray[82][186], dotarray[83][186], dotarray[84][186], dotarray[85][186], dotarray[86][186], dotarray[87][186], dotarray[88][186], dotarray[89][186], dotarray[90][186], dotarray[91][186], dotarray[92][186], dotarray[93][186], dotarray[94][186], dotarray[95][186], dotarray[96][186], dotarray[97][186], dotarray[98][186], dotarray[99][186], dotarray[100][186], dotarray[101][186], dotarray[102][186], dotarray[103][186], dotarray[104][186], dotarray[105][186], dotarray[106][186], dotarray[107][186], dotarray[108][186], dotarray[109][186], dotarray[110][186], dotarray[111][186], dotarray[112][186], dotarray[113][186], dotarray[114][186], dotarray[115][186], dotarray[116][186], dotarray[117][186], dotarray[118][186], dotarray[119][186], dotarray[120][186], dotarray[121][186], dotarray[122][186], dotarray[123][186], dotarray[124][186], dotarray[125][186], dotarray[126][186], dotarray[127][186]};
assign dot_col_187 = {dotarray[0][187], dotarray[1][187], dotarray[2][187], dotarray[3][187], dotarray[4][187], dotarray[5][187], dotarray[6][187], dotarray[7][187], dotarray[8][187], dotarray[9][187], dotarray[10][187], dotarray[11][187], dotarray[12][187], dotarray[13][187], dotarray[14][187], dotarray[15][187], dotarray[16][187], dotarray[17][187], dotarray[18][187], dotarray[19][187], dotarray[20][187], dotarray[21][187], dotarray[22][187], dotarray[23][187], dotarray[24][187], dotarray[25][187], dotarray[26][187], dotarray[27][187], dotarray[28][187], dotarray[29][187], dotarray[30][187], dotarray[31][187], dotarray[32][187], dotarray[33][187], dotarray[34][187], dotarray[35][187], dotarray[36][187], dotarray[37][187], dotarray[38][187], dotarray[39][187], dotarray[40][187], dotarray[41][187], dotarray[42][187], dotarray[43][187], dotarray[44][187], dotarray[45][187], dotarray[46][187], dotarray[47][187], dotarray[48][187], dotarray[49][187], dotarray[50][187], dotarray[51][187], dotarray[52][187], dotarray[53][187], dotarray[54][187], dotarray[55][187], dotarray[56][187], dotarray[57][187], dotarray[58][187], dotarray[59][187], dotarray[60][187], dotarray[61][187], dotarray[62][187], dotarray[63][187], dotarray[64][187], dotarray[65][187], dotarray[66][187], dotarray[67][187], dotarray[68][187], dotarray[69][187], dotarray[70][187], dotarray[71][187], dotarray[72][187], dotarray[73][187], dotarray[74][187], dotarray[75][187], dotarray[76][187], dotarray[77][187], dotarray[78][187], dotarray[79][187], dotarray[80][187], dotarray[81][187], dotarray[82][187], dotarray[83][187], dotarray[84][187], dotarray[85][187], dotarray[86][187], dotarray[87][187], dotarray[88][187], dotarray[89][187], dotarray[90][187], dotarray[91][187], dotarray[92][187], dotarray[93][187], dotarray[94][187], dotarray[95][187], dotarray[96][187], dotarray[97][187], dotarray[98][187], dotarray[99][187], dotarray[100][187], dotarray[101][187], dotarray[102][187], dotarray[103][187], dotarray[104][187], dotarray[105][187], dotarray[106][187], dotarray[107][187], dotarray[108][187], dotarray[109][187], dotarray[110][187], dotarray[111][187], dotarray[112][187], dotarray[113][187], dotarray[114][187], dotarray[115][187], dotarray[116][187], dotarray[117][187], dotarray[118][187], dotarray[119][187], dotarray[120][187], dotarray[121][187], dotarray[122][187], dotarray[123][187], dotarray[124][187], dotarray[125][187], dotarray[126][187], dotarray[127][187]};
assign dot_col_188 = {dotarray[0][188], dotarray[1][188], dotarray[2][188], dotarray[3][188], dotarray[4][188], dotarray[5][188], dotarray[6][188], dotarray[7][188], dotarray[8][188], dotarray[9][188], dotarray[10][188], dotarray[11][188], dotarray[12][188], dotarray[13][188], dotarray[14][188], dotarray[15][188], dotarray[16][188], dotarray[17][188], dotarray[18][188], dotarray[19][188], dotarray[20][188], dotarray[21][188], dotarray[22][188], dotarray[23][188], dotarray[24][188], dotarray[25][188], dotarray[26][188], dotarray[27][188], dotarray[28][188], dotarray[29][188], dotarray[30][188], dotarray[31][188], dotarray[32][188], dotarray[33][188], dotarray[34][188], dotarray[35][188], dotarray[36][188], dotarray[37][188], dotarray[38][188], dotarray[39][188], dotarray[40][188], dotarray[41][188], dotarray[42][188], dotarray[43][188], dotarray[44][188], dotarray[45][188], dotarray[46][188], dotarray[47][188], dotarray[48][188], dotarray[49][188], dotarray[50][188], dotarray[51][188], dotarray[52][188], dotarray[53][188], dotarray[54][188], dotarray[55][188], dotarray[56][188], dotarray[57][188], dotarray[58][188], dotarray[59][188], dotarray[60][188], dotarray[61][188], dotarray[62][188], dotarray[63][188], dotarray[64][188], dotarray[65][188], dotarray[66][188], dotarray[67][188], dotarray[68][188], dotarray[69][188], dotarray[70][188], dotarray[71][188], dotarray[72][188], dotarray[73][188], dotarray[74][188], dotarray[75][188], dotarray[76][188], dotarray[77][188], dotarray[78][188], dotarray[79][188], dotarray[80][188], dotarray[81][188], dotarray[82][188], dotarray[83][188], dotarray[84][188], dotarray[85][188], dotarray[86][188], dotarray[87][188], dotarray[88][188], dotarray[89][188], dotarray[90][188], dotarray[91][188], dotarray[92][188], dotarray[93][188], dotarray[94][188], dotarray[95][188], dotarray[96][188], dotarray[97][188], dotarray[98][188], dotarray[99][188], dotarray[100][188], dotarray[101][188], dotarray[102][188], dotarray[103][188], dotarray[104][188], dotarray[105][188], dotarray[106][188], dotarray[107][188], dotarray[108][188], dotarray[109][188], dotarray[110][188], dotarray[111][188], dotarray[112][188], dotarray[113][188], dotarray[114][188], dotarray[115][188], dotarray[116][188], dotarray[117][188], dotarray[118][188], dotarray[119][188], dotarray[120][188], dotarray[121][188], dotarray[122][188], dotarray[123][188], dotarray[124][188], dotarray[125][188], dotarray[126][188], dotarray[127][188]};
assign dot_col_189 = {dotarray[0][189], dotarray[1][189], dotarray[2][189], dotarray[3][189], dotarray[4][189], dotarray[5][189], dotarray[6][189], dotarray[7][189], dotarray[8][189], dotarray[9][189], dotarray[10][189], dotarray[11][189], dotarray[12][189], dotarray[13][189], dotarray[14][189], dotarray[15][189], dotarray[16][189], dotarray[17][189], dotarray[18][189], dotarray[19][189], dotarray[20][189], dotarray[21][189], dotarray[22][189], dotarray[23][189], dotarray[24][189], dotarray[25][189], dotarray[26][189], dotarray[27][189], dotarray[28][189], dotarray[29][189], dotarray[30][189], dotarray[31][189], dotarray[32][189], dotarray[33][189], dotarray[34][189], dotarray[35][189], dotarray[36][189], dotarray[37][189], dotarray[38][189], dotarray[39][189], dotarray[40][189], dotarray[41][189], dotarray[42][189], dotarray[43][189], dotarray[44][189], dotarray[45][189], dotarray[46][189], dotarray[47][189], dotarray[48][189], dotarray[49][189], dotarray[50][189], dotarray[51][189], dotarray[52][189], dotarray[53][189], dotarray[54][189], dotarray[55][189], dotarray[56][189], dotarray[57][189], dotarray[58][189], dotarray[59][189], dotarray[60][189], dotarray[61][189], dotarray[62][189], dotarray[63][189], dotarray[64][189], dotarray[65][189], dotarray[66][189], dotarray[67][189], dotarray[68][189], dotarray[69][189], dotarray[70][189], dotarray[71][189], dotarray[72][189], dotarray[73][189], dotarray[74][189], dotarray[75][189], dotarray[76][189], dotarray[77][189], dotarray[78][189], dotarray[79][189], dotarray[80][189], dotarray[81][189], dotarray[82][189], dotarray[83][189], dotarray[84][189], dotarray[85][189], dotarray[86][189], dotarray[87][189], dotarray[88][189], dotarray[89][189], dotarray[90][189], dotarray[91][189], dotarray[92][189], dotarray[93][189], dotarray[94][189], dotarray[95][189], dotarray[96][189], dotarray[97][189], dotarray[98][189], dotarray[99][189], dotarray[100][189], dotarray[101][189], dotarray[102][189], dotarray[103][189], dotarray[104][189], dotarray[105][189], dotarray[106][189], dotarray[107][189], dotarray[108][189], dotarray[109][189], dotarray[110][189], dotarray[111][189], dotarray[112][189], dotarray[113][189], dotarray[114][189], dotarray[115][189], dotarray[116][189], dotarray[117][189], dotarray[118][189], dotarray[119][189], dotarray[120][189], dotarray[121][189], dotarray[122][189], dotarray[123][189], dotarray[124][189], dotarray[125][189], dotarray[126][189], dotarray[127][189]};
assign dot_col_190 = {dotarray[0][190], dotarray[1][190], dotarray[2][190], dotarray[3][190], dotarray[4][190], dotarray[5][190], dotarray[6][190], dotarray[7][190], dotarray[8][190], dotarray[9][190], dotarray[10][190], dotarray[11][190], dotarray[12][190], dotarray[13][190], dotarray[14][190], dotarray[15][190], dotarray[16][190], dotarray[17][190], dotarray[18][190], dotarray[19][190], dotarray[20][190], dotarray[21][190], dotarray[22][190], dotarray[23][190], dotarray[24][190], dotarray[25][190], dotarray[26][190], dotarray[27][190], dotarray[28][190], dotarray[29][190], dotarray[30][190], dotarray[31][190], dotarray[32][190], dotarray[33][190], dotarray[34][190], dotarray[35][190], dotarray[36][190], dotarray[37][190], dotarray[38][190], dotarray[39][190], dotarray[40][190], dotarray[41][190], dotarray[42][190], dotarray[43][190], dotarray[44][190], dotarray[45][190], dotarray[46][190], dotarray[47][190], dotarray[48][190], dotarray[49][190], dotarray[50][190], dotarray[51][190], dotarray[52][190], dotarray[53][190], dotarray[54][190], dotarray[55][190], dotarray[56][190], dotarray[57][190], dotarray[58][190], dotarray[59][190], dotarray[60][190], dotarray[61][190], dotarray[62][190], dotarray[63][190], dotarray[64][190], dotarray[65][190], dotarray[66][190], dotarray[67][190], dotarray[68][190], dotarray[69][190], dotarray[70][190], dotarray[71][190], dotarray[72][190], dotarray[73][190], dotarray[74][190], dotarray[75][190], dotarray[76][190], dotarray[77][190], dotarray[78][190], dotarray[79][190], dotarray[80][190], dotarray[81][190], dotarray[82][190], dotarray[83][190], dotarray[84][190], dotarray[85][190], dotarray[86][190], dotarray[87][190], dotarray[88][190], dotarray[89][190], dotarray[90][190], dotarray[91][190], dotarray[92][190], dotarray[93][190], dotarray[94][190], dotarray[95][190], dotarray[96][190], dotarray[97][190], dotarray[98][190], dotarray[99][190], dotarray[100][190], dotarray[101][190], dotarray[102][190], dotarray[103][190], dotarray[104][190], dotarray[105][190], dotarray[106][190], dotarray[107][190], dotarray[108][190], dotarray[109][190], dotarray[110][190], dotarray[111][190], dotarray[112][190], dotarray[113][190], dotarray[114][190], dotarray[115][190], dotarray[116][190], dotarray[117][190], dotarray[118][190], dotarray[119][190], dotarray[120][190], dotarray[121][190], dotarray[122][190], dotarray[123][190], dotarray[124][190], dotarray[125][190], dotarray[126][190], dotarray[127][190]};
assign dot_col_191 = {dotarray[0][191], dotarray[1][191], dotarray[2][191], dotarray[3][191], dotarray[4][191], dotarray[5][191], dotarray[6][191], dotarray[7][191], dotarray[8][191], dotarray[9][191], dotarray[10][191], dotarray[11][191], dotarray[12][191], dotarray[13][191], dotarray[14][191], dotarray[15][191], dotarray[16][191], dotarray[17][191], dotarray[18][191], dotarray[19][191], dotarray[20][191], dotarray[21][191], dotarray[22][191], dotarray[23][191], dotarray[24][191], dotarray[25][191], dotarray[26][191], dotarray[27][191], dotarray[28][191], dotarray[29][191], dotarray[30][191], dotarray[31][191], dotarray[32][191], dotarray[33][191], dotarray[34][191], dotarray[35][191], dotarray[36][191], dotarray[37][191], dotarray[38][191], dotarray[39][191], dotarray[40][191], dotarray[41][191], dotarray[42][191], dotarray[43][191], dotarray[44][191], dotarray[45][191], dotarray[46][191], dotarray[47][191], dotarray[48][191], dotarray[49][191], dotarray[50][191], dotarray[51][191], dotarray[52][191], dotarray[53][191], dotarray[54][191], dotarray[55][191], dotarray[56][191], dotarray[57][191], dotarray[58][191], dotarray[59][191], dotarray[60][191], dotarray[61][191], dotarray[62][191], dotarray[63][191], dotarray[64][191], dotarray[65][191], dotarray[66][191], dotarray[67][191], dotarray[68][191], dotarray[69][191], dotarray[70][191], dotarray[71][191], dotarray[72][191], dotarray[73][191], dotarray[74][191], dotarray[75][191], dotarray[76][191], dotarray[77][191], dotarray[78][191], dotarray[79][191], dotarray[80][191], dotarray[81][191], dotarray[82][191], dotarray[83][191], dotarray[84][191], dotarray[85][191], dotarray[86][191], dotarray[87][191], dotarray[88][191], dotarray[89][191], dotarray[90][191], dotarray[91][191], dotarray[92][191], dotarray[93][191], dotarray[94][191], dotarray[95][191], dotarray[96][191], dotarray[97][191], dotarray[98][191], dotarray[99][191], dotarray[100][191], dotarray[101][191], dotarray[102][191], dotarray[103][191], dotarray[104][191], dotarray[105][191], dotarray[106][191], dotarray[107][191], dotarray[108][191], dotarray[109][191], dotarray[110][191], dotarray[111][191], dotarray[112][191], dotarray[113][191], dotarray[114][191], dotarray[115][191], dotarray[116][191], dotarray[117][191], dotarray[118][191], dotarray[119][191], dotarray[120][191], dotarray[121][191], dotarray[122][191], dotarray[123][191], dotarray[124][191], dotarray[125][191], dotarray[126][191], dotarray[127][191]};
assign dot_col_192 = {dotarray[0][192], dotarray[1][192], dotarray[2][192], dotarray[3][192], dotarray[4][192], dotarray[5][192], dotarray[6][192], dotarray[7][192], dotarray[8][192], dotarray[9][192], dotarray[10][192], dotarray[11][192], dotarray[12][192], dotarray[13][192], dotarray[14][192], dotarray[15][192], dotarray[16][192], dotarray[17][192], dotarray[18][192], dotarray[19][192], dotarray[20][192], dotarray[21][192], dotarray[22][192], dotarray[23][192], dotarray[24][192], dotarray[25][192], dotarray[26][192], dotarray[27][192], dotarray[28][192], dotarray[29][192], dotarray[30][192], dotarray[31][192], dotarray[32][192], dotarray[33][192], dotarray[34][192], dotarray[35][192], dotarray[36][192], dotarray[37][192], dotarray[38][192], dotarray[39][192], dotarray[40][192], dotarray[41][192], dotarray[42][192], dotarray[43][192], dotarray[44][192], dotarray[45][192], dotarray[46][192], dotarray[47][192], dotarray[48][192], dotarray[49][192], dotarray[50][192], dotarray[51][192], dotarray[52][192], dotarray[53][192], dotarray[54][192], dotarray[55][192], dotarray[56][192], dotarray[57][192], dotarray[58][192], dotarray[59][192], dotarray[60][192], dotarray[61][192], dotarray[62][192], dotarray[63][192], dotarray[64][192], dotarray[65][192], dotarray[66][192], dotarray[67][192], dotarray[68][192], dotarray[69][192], dotarray[70][192], dotarray[71][192], dotarray[72][192], dotarray[73][192], dotarray[74][192], dotarray[75][192], dotarray[76][192], dotarray[77][192], dotarray[78][192], dotarray[79][192], dotarray[80][192], dotarray[81][192], dotarray[82][192], dotarray[83][192], dotarray[84][192], dotarray[85][192], dotarray[86][192], dotarray[87][192], dotarray[88][192], dotarray[89][192], dotarray[90][192], dotarray[91][192], dotarray[92][192], dotarray[93][192], dotarray[94][192], dotarray[95][192], dotarray[96][192], dotarray[97][192], dotarray[98][192], dotarray[99][192], dotarray[100][192], dotarray[101][192], dotarray[102][192], dotarray[103][192], dotarray[104][192], dotarray[105][192], dotarray[106][192], dotarray[107][192], dotarray[108][192], dotarray[109][192], dotarray[110][192], dotarray[111][192], dotarray[112][192], dotarray[113][192], dotarray[114][192], dotarray[115][192], dotarray[116][192], dotarray[117][192], dotarray[118][192], dotarray[119][192], dotarray[120][192], dotarray[121][192], dotarray[122][192], dotarray[123][192], dotarray[124][192], dotarray[125][192], dotarray[126][192], dotarray[127][192]};
assign dot_col_193 = {dotarray[0][193], dotarray[1][193], dotarray[2][193], dotarray[3][193], dotarray[4][193], dotarray[5][193], dotarray[6][193], dotarray[7][193], dotarray[8][193], dotarray[9][193], dotarray[10][193], dotarray[11][193], dotarray[12][193], dotarray[13][193], dotarray[14][193], dotarray[15][193], dotarray[16][193], dotarray[17][193], dotarray[18][193], dotarray[19][193], dotarray[20][193], dotarray[21][193], dotarray[22][193], dotarray[23][193], dotarray[24][193], dotarray[25][193], dotarray[26][193], dotarray[27][193], dotarray[28][193], dotarray[29][193], dotarray[30][193], dotarray[31][193], dotarray[32][193], dotarray[33][193], dotarray[34][193], dotarray[35][193], dotarray[36][193], dotarray[37][193], dotarray[38][193], dotarray[39][193], dotarray[40][193], dotarray[41][193], dotarray[42][193], dotarray[43][193], dotarray[44][193], dotarray[45][193], dotarray[46][193], dotarray[47][193], dotarray[48][193], dotarray[49][193], dotarray[50][193], dotarray[51][193], dotarray[52][193], dotarray[53][193], dotarray[54][193], dotarray[55][193], dotarray[56][193], dotarray[57][193], dotarray[58][193], dotarray[59][193], dotarray[60][193], dotarray[61][193], dotarray[62][193], dotarray[63][193], dotarray[64][193], dotarray[65][193], dotarray[66][193], dotarray[67][193], dotarray[68][193], dotarray[69][193], dotarray[70][193], dotarray[71][193], dotarray[72][193], dotarray[73][193], dotarray[74][193], dotarray[75][193], dotarray[76][193], dotarray[77][193], dotarray[78][193], dotarray[79][193], dotarray[80][193], dotarray[81][193], dotarray[82][193], dotarray[83][193], dotarray[84][193], dotarray[85][193], dotarray[86][193], dotarray[87][193], dotarray[88][193], dotarray[89][193], dotarray[90][193], dotarray[91][193], dotarray[92][193], dotarray[93][193], dotarray[94][193], dotarray[95][193], dotarray[96][193], dotarray[97][193], dotarray[98][193], dotarray[99][193], dotarray[100][193], dotarray[101][193], dotarray[102][193], dotarray[103][193], dotarray[104][193], dotarray[105][193], dotarray[106][193], dotarray[107][193], dotarray[108][193], dotarray[109][193], dotarray[110][193], dotarray[111][193], dotarray[112][193], dotarray[113][193], dotarray[114][193], dotarray[115][193], dotarray[116][193], dotarray[117][193], dotarray[118][193], dotarray[119][193], dotarray[120][193], dotarray[121][193], dotarray[122][193], dotarray[123][193], dotarray[124][193], dotarray[125][193], dotarray[126][193], dotarray[127][193]};
assign dot_col_194 = {dotarray[0][194], dotarray[1][194], dotarray[2][194], dotarray[3][194], dotarray[4][194], dotarray[5][194], dotarray[6][194], dotarray[7][194], dotarray[8][194], dotarray[9][194], dotarray[10][194], dotarray[11][194], dotarray[12][194], dotarray[13][194], dotarray[14][194], dotarray[15][194], dotarray[16][194], dotarray[17][194], dotarray[18][194], dotarray[19][194], dotarray[20][194], dotarray[21][194], dotarray[22][194], dotarray[23][194], dotarray[24][194], dotarray[25][194], dotarray[26][194], dotarray[27][194], dotarray[28][194], dotarray[29][194], dotarray[30][194], dotarray[31][194], dotarray[32][194], dotarray[33][194], dotarray[34][194], dotarray[35][194], dotarray[36][194], dotarray[37][194], dotarray[38][194], dotarray[39][194], dotarray[40][194], dotarray[41][194], dotarray[42][194], dotarray[43][194], dotarray[44][194], dotarray[45][194], dotarray[46][194], dotarray[47][194], dotarray[48][194], dotarray[49][194], dotarray[50][194], dotarray[51][194], dotarray[52][194], dotarray[53][194], dotarray[54][194], dotarray[55][194], dotarray[56][194], dotarray[57][194], dotarray[58][194], dotarray[59][194], dotarray[60][194], dotarray[61][194], dotarray[62][194], dotarray[63][194], dotarray[64][194], dotarray[65][194], dotarray[66][194], dotarray[67][194], dotarray[68][194], dotarray[69][194], dotarray[70][194], dotarray[71][194], dotarray[72][194], dotarray[73][194], dotarray[74][194], dotarray[75][194], dotarray[76][194], dotarray[77][194], dotarray[78][194], dotarray[79][194], dotarray[80][194], dotarray[81][194], dotarray[82][194], dotarray[83][194], dotarray[84][194], dotarray[85][194], dotarray[86][194], dotarray[87][194], dotarray[88][194], dotarray[89][194], dotarray[90][194], dotarray[91][194], dotarray[92][194], dotarray[93][194], dotarray[94][194], dotarray[95][194], dotarray[96][194], dotarray[97][194], dotarray[98][194], dotarray[99][194], dotarray[100][194], dotarray[101][194], dotarray[102][194], dotarray[103][194], dotarray[104][194], dotarray[105][194], dotarray[106][194], dotarray[107][194], dotarray[108][194], dotarray[109][194], dotarray[110][194], dotarray[111][194], dotarray[112][194], dotarray[113][194], dotarray[114][194], dotarray[115][194], dotarray[116][194], dotarray[117][194], dotarray[118][194], dotarray[119][194], dotarray[120][194], dotarray[121][194], dotarray[122][194], dotarray[123][194], dotarray[124][194], dotarray[125][194], dotarray[126][194], dotarray[127][194]};
assign dot_col_195 = {dotarray[0][195], dotarray[1][195], dotarray[2][195], dotarray[3][195], dotarray[4][195], dotarray[5][195], dotarray[6][195], dotarray[7][195], dotarray[8][195], dotarray[9][195], dotarray[10][195], dotarray[11][195], dotarray[12][195], dotarray[13][195], dotarray[14][195], dotarray[15][195], dotarray[16][195], dotarray[17][195], dotarray[18][195], dotarray[19][195], dotarray[20][195], dotarray[21][195], dotarray[22][195], dotarray[23][195], dotarray[24][195], dotarray[25][195], dotarray[26][195], dotarray[27][195], dotarray[28][195], dotarray[29][195], dotarray[30][195], dotarray[31][195], dotarray[32][195], dotarray[33][195], dotarray[34][195], dotarray[35][195], dotarray[36][195], dotarray[37][195], dotarray[38][195], dotarray[39][195], dotarray[40][195], dotarray[41][195], dotarray[42][195], dotarray[43][195], dotarray[44][195], dotarray[45][195], dotarray[46][195], dotarray[47][195], dotarray[48][195], dotarray[49][195], dotarray[50][195], dotarray[51][195], dotarray[52][195], dotarray[53][195], dotarray[54][195], dotarray[55][195], dotarray[56][195], dotarray[57][195], dotarray[58][195], dotarray[59][195], dotarray[60][195], dotarray[61][195], dotarray[62][195], dotarray[63][195], dotarray[64][195], dotarray[65][195], dotarray[66][195], dotarray[67][195], dotarray[68][195], dotarray[69][195], dotarray[70][195], dotarray[71][195], dotarray[72][195], dotarray[73][195], dotarray[74][195], dotarray[75][195], dotarray[76][195], dotarray[77][195], dotarray[78][195], dotarray[79][195], dotarray[80][195], dotarray[81][195], dotarray[82][195], dotarray[83][195], dotarray[84][195], dotarray[85][195], dotarray[86][195], dotarray[87][195], dotarray[88][195], dotarray[89][195], dotarray[90][195], dotarray[91][195], dotarray[92][195], dotarray[93][195], dotarray[94][195], dotarray[95][195], dotarray[96][195], dotarray[97][195], dotarray[98][195], dotarray[99][195], dotarray[100][195], dotarray[101][195], dotarray[102][195], dotarray[103][195], dotarray[104][195], dotarray[105][195], dotarray[106][195], dotarray[107][195], dotarray[108][195], dotarray[109][195], dotarray[110][195], dotarray[111][195], dotarray[112][195], dotarray[113][195], dotarray[114][195], dotarray[115][195], dotarray[116][195], dotarray[117][195], dotarray[118][195], dotarray[119][195], dotarray[120][195], dotarray[121][195], dotarray[122][195], dotarray[123][195], dotarray[124][195], dotarray[125][195], dotarray[126][195], dotarray[127][195]};
assign dot_col_196 = {dotarray[0][196], dotarray[1][196], dotarray[2][196], dotarray[3][196], dotarray[4][196], dotarray[5][196], dotarray[6][196], dotarray[7][196], dotarray[8][196], dotarray[9][196], dotarray[10][196], dotarray[11][196], dotarray[12][196], dotarray[13][196], dotarray[14][196], dotarray[15][196], dotarray[16][196], dotarray[17][196], dotarray[18][196], dotarray[19][196], dotarray[20][196], dotarray[21][196], dotarray[22][196], dotarray[23][196], dotarray[24][196], dotarray[25][196], dotarray[26][196], dotarray[27][196], dotarray[28][196], dotarray[29][196], dotarray[30][196], dotarray[31][196], dotarray[32][196], dotarray[33][196], dotarray[34][196], dotarray[35][196], dotarray[36][196], dotarray[37][196], dotarray[38][196], dotarray[39][196], dotarray[40][196], dotarray[41][196], dotarray[42][196], dotarray[43][196], dotarray[44][196], dotarray[45][196], dotarray[46][196], dotarray[47][196], dotarray[48][196], dotarray[49][196], dotarray[50][196], dotarray[51][196], dotarray[52][196], dotarray[53][196], dotarray[54][196], dotarray[55][196], dotarray[56][196], dotarray[57][196], dotarray[58][196], dotarray[59][196], dotarray[60][196], dotarray[61][196], dotarray[62][196], dotarray[63][196], dotarray[64][196], dotarray[65][196], dotarray[66][196], dotarray[67][196], dotarray[68][196], dotarray[69][196], dotarray[70][196], dotarray[71][196], dotarray[72][196], dotarray[73][196], dotarray[74][196], dotarray[75][196], dotarray[76][196], dotarray[77][196], dotarray[78][196], dotarray[79][196], dotarray[80][196], dotarray[81][196], dotarray[82][196], dotarray[83][196], dotarray[84][196], dotarray[85][196], dotarray[86][196], dotarray[87][196], dotarray[88][196], dotarray[89][196], dotarray[90][196], dotarray[91][196], dotarray[92][196], dotarray[93][196], dotarray[94][196], dotarray[95][196], dotarray[96][196], dotarray[97][196], dotarray[98][196], dotarray[99][196], dotarray[100][196], dotarray[101][196], dotarray[102][196], dotarray[103][196], dotarray[104][196], dotarray[105][196], dotarray[106][196], dotarray[107][196], dotarray[108][196], dotarray[109][196], dotarray[110][196], dotarray[111][196], dotarray[112][196], dotarray[113][196], dotarray[114][196], dotarray[115][196], dotarray[116][196], dotarray[117][196], dotarray[118][196], dotarray[119][196], dotarray[120][196], dotarray[121][196], dotarray[122][196], dotarray[123][196], dotarray[124][196], dotarray[125][196], dotarray[126][196], dotarray[127][196]};
assign dot_col_197 = {dotarray[0][197], dotarray[1][197], dotarray[2][197], dotarray[3][197], dotarray[4][197], dotarray[5][197], dotarray[6][197], dotarray[7][197], dotarray[8][197], dotarray[9][197], dotarray[10][197], dotarray[11][197], dotarray[12][197], dotarray[13][197], dotarray[14][197], dotarray[15][197], dotarray[16][197], dotarray[17][197], dotarray[18][197], dotarray[19][197], dotarray[20][197], dotarray[21][197], dotarray[22][197], dotarray[23][197], dotarray[24][197], dotarray[25][197], dotarray[26][197], dotarray[27][197], dotarray[28][197], dotarray[29][197], dotarray[30][197], dotarray[31][197], dotarray[32][197], dotarray[33][197], dotarray[34][197], dotarray[35][197], dotarray[36][197], dotarray[37][197], dotarray[38][197], dotarray[39][197], dotarray[40][197], dotarray[41][197], dotarray[42][197], dotarray[43][197], dotarray[44][197], dotarray[45][197], dotarray[46][197], dotarray[47][197], dotarray[48][197], dotarray[49][197], dotarray[50][197], dotarray[51][197], dotarray[52][197], dotarray[53][197], dotarray[54][197], dotarray[55][197], dotarray[56][197], dotarray[57][197], dotarray[58][197], dotarray[59][197], dotarray[60][197], dotarray[61][197], dotarray[62][197], dotarray[63][197], dotarray[64][197], dotarray[65][197], dotarray[66][197], dotarray[67][197], dotarray[68][197], dotarray[69][197], dotarray[70][197], dotarray[71][197], dotarray[72][197], dotarray[73][197], dotarray[74][197], dotarray[75][197], dotarray[76][197], dotarray[77][197], dotarray[78][197], dotarray[79][197], dotarray[80][197], dotarray[81][197], dotarray[82][197], dotarray[83][197], dotarray[84][197], dotarray[85][197], dotarray[86][197], dotarray[87][197], dotarray[88][197], dotarray[89][197], dotarray[90][197], dotarray[91][197], dotarray[92][197], dotarray[93][197], dotarray[94][197], dotarray[95][197], dotarray[96][197], dotarray[97][197], dotarray[98][197], dotarray[99][197], dotarray[100][197], dotarray[101][197], dotarray[102][197], dotarray[103][197], dotarray[104][197], dotarray[105][197], dotarray[106][197], dotarray[107][197], dotarray[108][197], dotarray[109][197], dotarray[110][197], dotarray[111][197], dotarray[112][197], dotarray[113][197], dotarray[114][197], dotarray[115][197], dotarray[116][197], dotarray[117][197], dotarray[118][197], dotarray[119][197], dotarray[120][197], dotarray[121][197], dotarray[122][197], dotarray[123][197], dotarray[124][197], dotarray[125][197], dotarray[126][197], dotarray[127][197]};
assign dot_col_198 = {dotarray[0][198], dotarray[1][198], dotarray[2][198], dotarray[3][198], dotarray[4][198], dotarray[5][198], dotarray[6][198], dotarray[7][198], dotarray[8][198], dotarray[9][198], dotarray[10][198], dotarray[11][198], dotarray[12][198], dotarray[13][198], dotarray[14][198], dotarray[15][198], dotarray[16][198], dotarray[17][198], dotarray[18][198], dotarray[19][198], dotarray[20][198], dotarray[21][198], dotarray[22][198], dotarray[23][198], dotarray[24][198], dotarray[25][198], dotarray[26][198], dotarray[27][198], dotarray[28][198], dotarray[29][198], dotarray[30][198], dotarray[31][198], dotarray[32][198], dotarray[33][198], dotarray[34][198], dotarray[35][198], dotarray[36][198], dotarray[37][198], dotarray[38][198], dotarray[39][198], dotarray[40][198], dotarray[41][198], dotarray[42][198], dotarray[43][198], dotarray[44][198], dotarray[45][198], dotarray[46][198], dotarray[47][198], dotarray[48][198], dotarray[49][198], dotarray[50][198], dotarray[51][198], dotarray[52][198], dotarray[53][198], dotarray[54][198], dotarray[55][198], dotarray[56][198], dotarray[57][198], dotarray[58][198], dotarray[59][198], dotarray[60][198], dotarray[61][198], dotarray[62][198], dotarray[63][198], dotarray[64][198], dotarray[65][198], dotarray[66][198], dotarray[67][198], dotarray[68][198], dotarray[69][198], dotarray[70][198], dotarray[71][198], dotarray[72][198], dotarray[73][198], dotarray[74][198], dotarray[75][198], dotarray[76][198], dotarray[77][198], dotarray[78][198], dotarray[79][198], dotarray[80][198], dotarray[81][198], dotarray[82][198], dotarray[83][198], dotarray[84][198], dotarray[85][198], dotarray[86][198], dotarray[87][198], dotarray[88][198], dotarray[89][198], dotarray[90][198], dotarray[91][198], dotarray[92][198], dotarray[93][198], dotarray[94][198], dotarray[95][198], dotarray[96][198], dotarray[97][198], dotarray[98][198], dotarray[99][198], dotarray[100][198], dotarray[101][198], dotarray[102][198], dotarray[103][198], dotarray[104][198], dotarray[105][198], dotarray[106][198], dotarray[107][198], dotarray[108][198], dotarray[109][198], dotarray[110][198], dotarray[111][198], dotarray[112][198], dotarray[113][198], dotarray[114][198], dotarray[115][198], dotarray[116][198], dotarray[117][198], dotarray[118][198], dotarray[119][198], dotarray[120][198], dotarray[121][198], dotarray[122][198], dotarray[123][198], dotarray[124][198], dotarray[125][198], dotarray[126][198], dotarray[127][198]};
assign dot_col_199 = {dotarray[0][199], dotarray[1][199], dotarray[2][199], dotarray[3][199], dotarray[4][199], dotarray[5][199], dotarray[6][199], dotarray[7][199], dotarray[8][199], dotarray[9][199], dotarray[10][199], dotarray[11][199], dotarray[12][199], dotarray[13][199], dotarray[14][199], dotarray[15][199], dotarray[16][199], dotarray[17][199], dotarray[18][199], dotarray[19][199], dotarray[20][199], dotarray[21][199], dotarray[22][199], dotarray[23][199], dotarray[24][199], dotarray[25][199], dotarray[26][199], dotarray[27][199], dotarray[28][199], dotarray[29][199], dotarray[30][199], dotarray[31][199], dotarray[32][199], dotarray[33][199], dotarray[34][199], dotarray[35][199], dotarray[36][199], dotarray[37][199], dotarray[38][199], dotarray[39][199], dotarray[40][199], dotarray[41][199], dotarray[42][199], dotarray[43][199], dotarray[44][199], dotarray[45][199], dotarray[46][199], dotarray[47][199], dotarray[48][199], dotarray[49][199], dotarray[50][199], dotarray[51][199], dotarray[52][199], dotarray[53][199], dotarray[54][199], dotarray[55][199], dotarray[56][199], dotarray[57][199], dotarray[58][199], dotarray[59][199], dotarray[60][199], dotarray[61][199], dotarray[62][199], dotarray[63][199], dotarray[64][199], dotarray[65][199], dotarray[66][199], dotarray[67][199], dotarray[68][199], dotarray[69][199], dotarray[70][199], dotarray[71][199], dotarray[72][199], dotarray[73][199], dotarray[74][199], dotarray[75][199], dotarray[76][199], dotarray[77][199], dotarray[78][199], dotarray[79][199], dotarray[80][199], dotarray[81][199], dotarray[82][199], dotarray[83][199], dotarray[84][199], dotarray[85][199], dotarray[86][199], dotarray[87][199], dotarray[88][199], dotarray[89][199], dotarray[90][199], dotarray[91][199], dotarray[92][199], dotarray[93][199], dotarray[94][199], dotarray[95][199], dotarray[96][199], dotarray[97][199], dotarray[98][199], dotarray[99][199], dotarray[100][199], dotarray[101][199], dotarray[102][199], dotarray[103][199], dotarray[104][199], dotarray[105][199], dotarray[106][199], dotarray[107][199], dotarray[108][199], dotarray[109][199], dotarray[110][199], dotarray[111][199], dotarray[112][199], dotarray[113][199], dotarray[114][199], dotarray[115][199], dotarray[116][199], dotarray[117][199], dotarray[118][199], dotarray[119][199], dotarray[120][199], dotarray[121][199], dotarray[122][199], dotarray[123][199], dotarray[124][199], dotarray[125][199], dotarray[126][199], dotarray[127][199]};
assign dot_col_200 = {dotarray[0][200], dotarray[1][200], dotarray[2][200], dotarray[3][200], dotarray[4][200], dotarray[5][200], dotarray[6][200], dotarray[7][200], dotarray[8][200], dotarray[9][200], dotarray[10][200], dotarray[11][200], dotarray[12][200], dotarray[13][200], dotarray[14][200], dotarray[15][200], dotarray[16][200], dotarray[17][200], dotarray[18][200], dotarray[19][200], dotarray[20][200], dotarray[21][200], dotarray[22][200], dotarray[23][200], dotarray[24][200], dotarray[25][200], dotarray[26][200], dotarray[27][200], dotarray[28][200], dotarray[29][200], dotarray[30][200], dotarray[31][200], dotarray[32][200], dotarray[33][200], dotarray[34][200], dotarray[35][200], dotarray[36][200], dotarray[37][200], dotarray[38][200], dotarray[39][200], dotarray[40][200], dotarray[41][200], dotarray[42][200], dotarray[43][200], dotarray[44][200], dotarray[45][200], dotarray[46][200], dotarray[47][200], dotarray[48][200], dotarray[49][200], dotarray[50][200], dotarray[51][200], dotarray[52][200], dotarray[53][200], dotarray[54][200], dotarray[55][200], dotarray[56][200], dotarray[57][200], dotarray[58][200], dotarray[59][200], dotarray[60][200], dotarray[61][200], dotarray[62][200], dotarray[63][200], dotarray[64][200], dotarray[65][200], dotarray[66][200], dotarray[67][200], dotarray[68][200], dotarray[69][200], dotarray[70][200], dotarray[71][200], dotarray[72][200], dotarray[73][200], dotarray[74][200], dotarray[75][200], dotarray[76][200], dotarray[77][200], dotarray[78][200], dotarray[79][200], dotarray[80][200], dotarray[81][200], dotarray[82][200], dotarray[83][200], dotarray[84][200], dotarray[85][200], dotarray[86][200], dotarray[87][200], dotarray[88][200], dotarray[89][200], dotarray[90][200], dotarray[91][200], dotarray[92][200], dotarray[93][200], dotarray[94][200], dotarray[95][200], dotarray[96][200], dotarray[97][200], dotarray[98][200], dotarray[99][200], dotarray[100][200], dotarray[101][200], dotarray[102][200], dotarray[103][200], dotarray[104][200], dotarray[105][200], dotarray[106][200], dotarray[107][200], dotarray[108][200], dotarray[109][200], dotarray[110][200], dotarray[111][200], dotarray[112][200], dotarray[113][200], dotarray[114][200], dotarray[115][200], dotarray[116][200], dotarray[117][200], dotarray[118][200], dotarray[119][200], dotarray[120][200], dotarray[121][200], dotarray[122][200], dotarray[123][200], dotarray[124][200], dotarray[125][200], dotarray[126][200], dotarray[127][200]};
assign dot_col_201 = {dotarray[0][201], dotarray[1][201], dotarray[2][201], dotarray[3][201], dotarray[4][201], dotarray[5][201], dotarray[6][201], dotarray[7][201], dotarray[8][201], dotarray[9][201], dotarray[10][201], dotarray[11][201], dotarray[12][201], dotarray[13][201], dotarray[14][201], dotarray[15][201], dotarray[16][201], dotarray[17][201], dotarray[18][201], dotarray[19][201], dotarray[20][201], dotarray[21][201], dotarray[22][201], dotarray[23][201], dotarray[24][201], dotarray[25][201], dotarray[26][201], dotarray[27][201], dotarray[28][201], dotarray[29][201], dotarray[30][201], dotarray[31][201], dotarray[32][201], dotarray[33][201], dotarray[34][201], dotarray[35][201], dotarray[36][201], dotarray[37][201], dotarray[38][201], dotarray[39][201], dotarray[40][201], dotarray[41][201], dotarray[42][201], dotarray[43][201], dotarray[44][201], dotarray[45][201], dotarray[46][201], dotarray[47][201], dotarray[48][201], dotarray[49][201], dotarray[50][201], dotarray[51][201], dotarray[52][201], dotarray[53][201], dotarray[54][201], dotarray[55][201], dotarray[56][201], dotarray[57][201], dotarray[58][201], dotarray[59][201], dotarray[60][201], dotarray[61][201], dotarray[62][201], dotarray[63][201], dotarray[64][201], dotarray[65][201], dotarray[66][201], dotarray[67][201], dotarray[68][201], dotarray[69][201], dotarray[70][201], dotarray[71][201], dotarray[72][201], dotarray[73][201], dotarray[74][201], dotarray[75][201], dotarray[76][201], dotarray[77][201], dotarray[78][201], dotarray[79][201], dotarray[80][201], dotarray[81][201], dotarray[82][201], dotarray[83][201], dotarray[84][201], dotarray[85][201], dotarray[86][201], dotarray[87][201], dotarray[88][201], dotarray[89][201], dotarray[90][201], dotarray[91][201], dotarray[92][201], dotarray[93][201], dotarray[94][201], dotarray[95][201], dotarray[96][201], dotarray[97][201], dotarray[98][201], dotarray[99][201], dotarray[100][201], dotarray[101][201], dotarray[102][201], dotarray[103][201], dotarray[104][201], dotarray[105][201], dotarray[106][201], dotarray[107][201], dotarray[108][201], dotarray[109][201], dotarray[110][201], dotarray[111][201], dotarray[112][201], dotarray[113][201], dotarray[114][201], dotarray[115][201], dotarray[116][201], dotarray[117][201], dotarray[118][201], dotarray[119][201], dotarray[120][201], dotarray[121][201], dotarray[122][201], dotarray[123][201], dotarray[124][201], dotarray[125][201], dotarray[126][201], dotarray[127][201]};
assign dot_col_202 = {dotarray[0][202], dotarray[1][202], dotarray[2][202], dotarray[3][202], dotarray[4][202], dotarray[5][202], dotarray[6][202], dotarray[7][202], dotarray[8][202], dotarray[9][202], dotarray[10][202], dotarray[11][202], dotarray[12][202], dotarray[13][202], dotarray[14][202], dotarray[15][202], dotarray[16][202], dotarray[17][202], dotarray[18][202], dotarray[19][202], dotarray[20][202], dotarray[21][202], dotarray[22][202], dotarray[23][202], dotarray[24][202], dotarray[25][202], dotarray[26][202], dotarray[27][202], dotarray[28][202], dotarray[29][202], dotarray[30][202], dotarray[31][202], dotarray[32][202], dotarray[33][202], dotarray[34][202], dotarray[35][202], dotarray[36][202], dotarray[37][202], dotarray[38][202], dotarray[39][202], dotarray[40][202], dotarray[41][202], dotarray[42][202], dotarray[43][202], dotarray[44][202], dotarray[45][202], dotarray[46][202], dotarray[47][202], dotarray[48][202], dotarray[49][202], dotarray[50][202], dotarray[51][202], dotarray[52][202], dotarray[53][202], dotarray[54][202], dotarray[55][202], dotarray[56][202], dotarray[57][202], dotarray[58][202], dotarray[59][202], dotarray[60][202], dotarray[61][202], dotarray[62][202], dotarray[63][202], dotarray[64][202], dotarray[65][202], dotarray[66][202], dotarray[67][202], dotarray[68][202], dotarray[69][202], dotarray[70][202], dotarray[71][202], dotarray[72][202], dotarray[73][202], dotarray[74][202], dotarray[75][202], dotarray[76][202], dotarray[77][202], dotarray[78][202], dotarray[79][202], dotarray[80][202], dotarray[81][202], dotarray[82][202], dotarray[83][202], dotarray[84][202], dotarray[85][202], dotarray[86][202], dotarray[87][202], dotarray[88][202], dotarray[89][202], dotarray[90][202], dotarray[91][202], dotarray[92][202], dotarray[93][202], dotarray[94][202], dotarray[95][202], dotarray[96][202], dotarray[97][202], dotarray[98][202], dotarray[99][202], dotarray[100][202], dotarray[101][202], dotarray[102][202], dotarray[103][202], dotarray[104][202], dotarray[105][202], dotarray[106][202], dotarray[107][202], dotarray[108][202], dotarray[109][202], dotarray[110][202], dotarray[111][202], dotarray[112][202], dotarray[113][202], dotarray[114][202], dotarray[115][202], dotarray[116][202], dotarray[117][202], dotarray[118][202], dotarray[119][202], dotarray[120][202], dotarray[121][202], dotarray[122][202], dotarray[123][202], dotarray[124][202], dotarray[125][202], dotarray[126][202], dotarray[127][202]};
assign dot_col_203 = {dotarray[0][203], dotarray[1][203], dotarray[2][203], dotarray[3][203], dotarray[4][203], dotarray[5][203], dotarray[6][203], dotarray[7][203], dotarray[8][203], dotarray[9][203], dotarray[10][203], dotarray[11][203], dotarray[12][203], dotarray[13][203], dotarray[14][203], dotarray[15][203], dotarray[16][203], dotarray[17][203], dotarray[18][203], dotarray[19][203], dotarray[20][203], dotarray[21][203], dotarray[22][203], dotarray[23][203], dotarray[24][203], dotarray[25][203], dotarray[26][203], dotarray[27][203], dotarray[28][203], dotarray[29][203], dotarray[30][203], dotarray[31][203], dotarray[32][203], dotarray[33][203], dotarray[34][203], dotarray[35][203], dotarray[36][203], dotarray[37][203], dotarray[38][203], dotarray[39][203], dotarray[40][203], dotarray[41][203], dotarray[42][203], dotarray[43][203], dotarray[44][203], dotarray[45][203], dotarray[46][203], dotarray[47][203], dotarray[48][203], dotarray[49][203], dotarray[50][203], dotarray[51][203], dotarray[52][203], dotarray[53][203], dotarray[54][203], dotarray[55][203], dotarray[56][203], dotarray[57][203], dotarray[58][203], dotarray[59][203], dotarray[60][203], dotarray[61][203], dotarray[62][203], dotarray[63][203], dotarray[64][203], dotarray[65][203], dotarray[66][203], dotarray[67][203], dotarray[68][203], dotarray[69][203], dotarray[70][203], dotarray[71][203], dotarray[72][203], dotarray[73][203], dotarray[74][203], dotarray[75][203], dotarray[76][203], dotarray[77][203], dotarray[78][203], dotarray[79][203], dotarray[80][203], dotarray[81][203], dotarray[82][203], dotarray[83][203], dotarray[84][203], dotarray[85][203], dotarray[86][203], dotarray[87][203], dotarray[88][203], dotarray[89][203], dotarray[90][203], dotarray[91][203], dotarray[92][203], dotarray[93][203], dotarray[94][203], dotarray[95][203], dotarray[96][203], dotarray[97][203], dotarray[98][203], dotarray[99][203], dotarray[100][203], dotarray[101][203], dotarray[102][203], dotarray[103][203], dotarray[104][203], dotarray[105][203], dotarray[106][203], dotarray[107][203], dotarray[108][203], dotarray[109][203], dotarray[110][203], dotarray[111][203], dotarray[112][203], dotarray[113][203], dotarray[114][203], dotarray[115][203], dotarray[116][203], dotarray[117][203], dotarray[118][203], dotarray[119][203], dotarray[120][203], dotarray[121][203], dotarray[122][203], dotarray[123][203], dotarray[124][203], dotarray[125][203], dotarray[126][203], dotarray[127][203]};
assign dot_col_204 = {dotarray[0][204], dotarray[1][204], dotarray[2][204], dotarray[3][204], dotarray[4][204], dotarray[5][204], dotarray[6][204], dotarray[7][204], dotarray[8][204], dotarray[9][204], dotarray[10][204], dotarray[11][204], dotarray[12][204], dotarray[13][204], dotarray[14][204], dotarray[15][204], dotarray[16][204], dotarray[17][204], dotarray[18][204], dotarray[19][204], dotarray[20][204], dotarray[21][204], dotarray[22][204], dotarray[23][204], dotarray[24][204], dotarray[25][204], dotarray[26][204], dotarray[27][204], dotarray[28][204], dotarray[29][204], dotarray[30][204], dotarray[31][204], dotarray[32][204], dotarray[33][204], dotarray[34][204], dotarray[35][204], dotarray[36][204], dotarray[37][204], dotarray[38][204], dotarray[39][204], dotarray[40][204], dotarray[41][204], dotarray[42][204], dotarray[43][204], dotarray[44][204], dotarray[45][204], dotarray[46][204], dotarray[47][204], dotarray[48][204], dotarray[49][204], dotarray[50][204], dotarray[51][204], dotarray[52][204], dotarray[53][204], dotarray[54][204], dotarray[55][204], dotarray[56][204], dotarray[57][204], dotarray[58][204], dotarray[59][204], dotarray[60][204], dotarray[61][204], dotarray[62][204], dotarray[63][204], dotarray[64][204], dotarray[65][204], dotarray[66][204], dotarray[67][204], dotarray[68][204], dotarray[69][204], dotarray[70][204], dotarray[71][204], dotarray[72][204], dotarray[73][204], dotarray[74][204], dotarray[75][204], dotarray[76][204], dotarray[77][204], dotarray[78][204], dotarray[79][204], dotarray[80][204], dotarray[81][204], dotarray[82][204], dotarray[83][204], dotarray[84][204], dotarray[85][204], dotarray[86][204], dotarray[87][204], dotarray[88][204], dotarray[89][204], dotarray[90][204], dotarray[91][204], dotarray[92][204], dotarray[93][204], dotarray[94][204], dotarray[95][204], dotarray[96][204], dotarray[97][204], dotarray[98][204], dotarray[99][204], dotarray[100][204], dotarray[101][204], dotarray[102][204], dotarray[103][204], dotarray[104][204], dotarray[105][204], dotarray[106][204], dotarray[107][204], dotarray[108][204], dotarray[109][204], dotarray[110][204], dotarray[111][204], dotarray[112][204], dotarray[113][204], dotarray[114][204], dotarray[115][204], dotarray[116][204], dotarray[117][204], dotarray[118][204], dotarray[119][204], dotarray[120][204], dotarray[121][204], dotarray[122][204], dotarray[123][204], dotarray[124][204], dotarray[125][204], dotarray[126][204], dotarray[127][204]};
assign dot_col_205 = {dotarray[0][205], dotarray[1][205], dotarray[2][205], dotarray[3][205], dotarray[4][205], dotarray[5][205], dotarray[6][205], dotarray[7][205], dotarray[8][205], dotarray[9][205], dotarray[10][205], dotarray[11][205], dotarray[12][205], dotarray[13][205], dotarray[14][205], dotarray[15][205], dotarray[16][205], dotarray[17][205], dotarray[18][205], dotarray[19][205], dotarray[20][205], dotarray[21][205], dotarray[22][205], dotarray[23][205], dotarray[24][205], dotarray[25][205], dotarray[26][205], dotarray[27][205], dotarray[28][205], dotarray[29][205], dotarray[30][205], dotarray[31][205], dotarray[32][205], dotarray[33][205], dotarray[34][205], dotarray[35][205], dotarray[36][205], dotarray[37][205], dotarray[38][205], dotarray[39][205], dotarray[40][205], dotarray[41][205], dotarray[42][205], dotarray[43][205], dotarray[44][205], dotarray[45][205], dotarray[46][205], dotarray[47][205], dotarray[48][205], dotarray[49][205], dotarray[50][205], dotarray[51][205], dotarray[52][205], dotarray[53][205], dotarray[54][205], dotarray[55][205], dotarray[56][205], dotarray[57][205], dotarray[58][205], dotarray[59][205], dotarray[60][205], dotarray[61][205], dotarray[62][205], dotarray[63][205], dotarray[64][205], dotarray[65][205], dotarray[66][205], dotarray[67][205], dotarray[68][205], dotarray[69][205], dotarray[70][205], dotarray[71][205], dotarray[72][205], dotarray[73][205], dotarray[74][205], dotarray[75][205], dotarray[76][205], dotarray[77][205], dotarray[78][205], dotarray[79][205], dotarray[80][205], dotarray[81][205], dotarray[82][205], dotarray[83][205], dotarray[84][205], dotarray[85][205], dotarray[86][205], dotarray[87][205], dotarray[88][205], dotarray[89][205], dotarray[90][205], dotarray[91][205], dotarray[92][205], dotarray[93][205], dotarray[94][205], dotarray[95][205], dotarray[96][205], dotarray[97][205], dotarray[98][205], dotarray[99][205], dotarray[100][205], dotarray[101][205], dotarray[102][205], dotarray[103][205], dotarray[104][205], dotarray[105][205], dotarray[106][205], dotarray[107][205], dotarray[108][205], dotarray[109][205], dotarray[110][205], dotarray[111][205], dotarray[112][205], dotarray[113][205], dotarray[114][205], dotarray[115][205], dotarray[116][205], dotarray[117][205], dotarray[118][205], dotarray[119][205], dotarray[120][205], dotarray[121][205], dotarray[122][205], dotarray[123][205], dotarray[124][205], dotarray[125][205], dotarray[126][205], dotarray[127][205]};
assign dot_col_206 = {dotarray[0][206], dotarray[1][206], dotarray[2][206], dotarray[3][206], dotarray[4][206], dotarray[5][206], dotarray[6][206], dotarray[7][206], dotarray[8][206], dotarray[9][206], dotarray[10][206], dotarray[11][206], dotarray[12][206], dotarray[13][206], dotarray[14][206], dotarray[15][206], dotarray[16][206], dotarray[17][206], dotarray[18][206], dotarray[19][206], dotarray[20][206], dotarray[21][206], dotarray[22][206], dotarray[23][206], dotarray[24][206], dotarray[25][206], dotarray[26][206], dotarray[27][206], dotarray[28][206], dotarray[29][206], dotarray[30][206], dotarray[31][206], dotarray[32][206], dotarray[33][206], dotarray[34][206], dotarray[35][206], dotarray[36][206], dotarray[37][206], dotarray[38][206], dotarray[39][206], dotarray[40][206], dotarray[41][206], dotarray[42][206], dotarray[43][206], dotarray[44][206], dotarray[45][206], dotarray[46][206], dotarray[47][206], dotarray[48][206], dotarray[49][206], dotarray[50][206], dotarray[51][206], dotarray[52][206], dotarray[53][206], dotarray[54][206], dotarray[55][206], dotarray[56][206], dotarray[57][206], dotarray[58][206], dotarray[59][206], dotarray[60][206], dotarray[61][206], dotarray[62][206], dotarray[63][206], dotarray[64][206], dotarray[65][206], dotarray[66][206], dotarray[67][206], dotarray[68][206], dotarray[69][206], dotarray[70][206], dotarray[71][206], dotarray[72][206], dotarray[73][206], dotarray[74][206], dotarray[75][206], dotarray[76][206], dotarray[77][206], dotarray[78][206], dotarray[79][206], dotarray[80][206], dotarray[81][206], dotarray[82][206], dotarray[83][206], dotarray[84][206], dotarray[85][206], dotarray[86][206], dotarray[87][206], dotarray[88][206], dotarray[89][206], dotarray[90][206], dotarray[91][206], dotarray[92][206], dotarray[93][206], dotarray[94][206], dotarray[95][206], dotarray[96][206], dotarray[97][206], dotarray[98][206], dotarray[99][206], dotarray[100][206], dotarray[101][206], dotarray[102][206], dotarray[103][206], dotarray[104][206], dotarray[105][206], dotarray[106][206], dotarray[107][206], dotarray[108][206], dotarray[109][206], dotarray[110][206], dotarray[111][206], dotarray[112][206], dotarray[113][206], dotarray[114][206], dotarray[115][206], dotarray[116][206], dotarray[117][206], dotarray[118][206], dotarray[119][206], dotarray[120][206], dotarray[121][206], dotarray[122][206], dotarray[123][206], dotarray[124][206], dotarray[125][206], dotarray[126][206], dotarray[127][206]};
assign dot_col_207 = {dotarray[0][207], dotarray[1][207], dotarray[2][207], dotarray[3][207], dotarray[4][207], dotarray[5][207], dotarray[6][207], dotarray[7][207], dotarray[8][207], dotarray[9][207], dotarray[10][207], dotarray[11][207], dotarray[12][207], dotarray[13][207], dotarray[14][207], dotarray[15][207], dotarray[16][207], dotarray[17][207], dotarray[18][207], dotarray[19][207], dotarray[20][207], dotarray[21][207], dotarray[22][207], dotarray[23][207], dotarray[24][207], dotarray[25][207], dotarray[26][207], dotarray[27][207], dotarray[28][207], dotarray[29][207], dotarray[30][207], dotarray[31][207], dotarray[32][207], dotarray[33][207], dotarray[34][207], dotarray[35][207], dotarray[36][207], dotarray[37][207], dotarray[38][207], dotarray[39][207], dotarray[40][207], dotarray[41][207], dotarray[42][207], dotarray[43][207], dotarray[44][207], dotarray[45][207], dotarray[46][207], dotarray[47][207], dotarray[48][207], dotarray[49][207], dotarray[50][207], dotarray[51][207], dotarray[52][207], dotarray[53][207], dotarray[54][207], dotarray[55][207], dotarray[56][207], dotarray[57][207], dotarray[58][207], dotarray[59][207], dotarray[60][207], dotarray[61][207], dotarray[62][207], dotarray[63][207], dotarray[64][207], dotarray[65][207], dotarray[66][207], dotarray[67][207], dotarray[68][207], dotarray[69][207], dotarray[70][207], dotarray[71][207], dotarray[72][207], dotarray[73][207], dotarray[74][207], dotarray[75][207], dotarray[76][207], dotarray[77][207], dotarray[78][207], dotarray[79][207], dotarray[80][207], dotarray[81][207], dotarray[82][207], dotarray[83][207], dotarray[84][207], dotarray[85][207], dotarray[86][207], dotarray[87][207], dotarray[88][207], dotarray[89][207], dotarray[90][207], dotarray[91][207], dotarray[92][207], dotarray[93][207], dotarray[94][207], dotarray[95][207], dotarray[96][207], dotarray[97][207], dotarray[98][207], dotarray[99][207], dotarray[100][207], dotarray[101][207], dotarray[102][207], dotarray[103][207], dotarray[104][207], dotarray[105][207], dotarray[106][207], dotarray[107][207], dotarray[108][207], dotarray[109][207], dotarray[110][207], dotarray[111][207], dotarray[112][207], dotarray[113][207], dotarray[114][207], dotarray[115][207], dotarray[116][207], dotarray[117][207], dotarray[118][207], dotarray[119][207], dotarray[120][207], dotarray[121][207], dotarray[122][207], dotarray[123][207], dotarray[124][207], dotarray[125][207], dotarray[126][207], dotarray[127][207]};
assign dot_col_208 = {dotarray[0][208], dotarray[1][208], dotarray[2][208], dotarray[3][208], dotarray[4][208], dotarray[5][208], dotarray[6][208], dotarray[7][208], dotarray[8][208], dotarray[9][208], dotarray[10][208], dotarray[11][208], dotarray[12][208], dotarray[13][208], dotarray[14][208], dotarray[15][208], dotarray[16][208], dotarray[17][208], dotarray[18][208], dotarray[19][208], dotarray[20][208], dotarray[21][208], dotarray[22][208], dotarray[23][208], dotarray[24][208], dotarray[25][208], dotarray[26][208], dotarray[27][208], dotarray[28][208], dotarray[29][208], dotarray[30][208], dotarray[31][208], dotarray[32][208], dotarray[33][208], dotarray[34][208], dotarray[35][208], dotarray[36][208], dotarray[37][208], dotarray[38][208], dotarray[39][208], dotarray[40][208], dotarray[41][208], dotarray[42][208], dotarray[43][208], dotarray[44][208], dotarray[45][208], dotarray[46][208], dotarray[47][208], dotarray[48][208], dotarray[49][208], dotarray[50][208], dotarray[51][208], dotarray[52][208], dotarray[53][208], dotarray[54][208], dotarray[55][208], dotarray[56][208], dotarray[57][208], dotarray[58][208], dotarray[59][208], dotarray[60][208], dotarray[61][208], dotarray[62][208], dotarray[63][208], dotarray[64][208], dotarray[65][208], dotarray[66][208], dotarray[67][208], dotarray[68][208], dotarray[69][208], dotarray[70][208], dotarray[71][208], dotarray[72][208], dotarray[73][208], dotarray[74][208], dotarray[75][208], dotarray[76][208], dotarray[77][208], dotarray[78][208], dotarray[79][208], dotarray[80][208], dotarray[81][208], dotarray[82][208], dotarray[83][208], dotarray[84][208], dotarray[85][208], dotarray[86][208], dotarray[87][208], dotarray[88][208], dotarray[89][208], dotarray[90][208], dotarray[91][208], dotarray[92][208], dotarray[93][208], dotarray[94][208], dotarray[95][208], dotarray[96][208], dotarray[97][208], dotarray[98][208], dotarray[99][208], dotarray[100][208], dotarray[101][208], dotarray[102][208], dotarray[103][208], dotarray[104][208], dotarray[105][208], dotarray[106][208], dotarray[107][208], dotarray[108][208], dotarray[109][208], dotarray[110][208], dotarray[111][208], dotarray[112][208], dotarray[113][208], dotarray[114][208], dotarray[115][208], dotarray[116][208], dotarray[117][208], dotarray[118][208], dotarray[119][208], dotarray[120][208], dotarray[121][208], dotarray[122][208], dotarray[123][208], dotarray[124][208], dotarray[125][208], dotarray[126][208], dotarray[127][208]};
assign dot_col_209 = {dotarray[0][209], dotarray[1][209], dotarray[2][209], dotarray[3][209], dotarray[4][209], dotarray[5][209], dotarray[6][209], dotarray[7][209], dotarray[8][209], dotarray[9][209], dotarray[10][209], dotarray[11][209], dotarray[12][209], dotarray[13][209], dotarray[14][209], dotarray[15][209], dotarray[16][209], dotarray[17][209], dotarray[18][209], dotarray[19][209], dotarray[20][209], dotarray[21][209], dotarray[22][209], dotarray[23][209], dotarray[24][209], dotarray[25][209], dotarray[26][209], dotarray[27][209], dotarray[28][209], dotarray[29][209], dotarray[30][209], dotarray[31][209], dotarray[32][209], dotarray[33][209], dotarray[34][209], dotarray[35][209], dotarray[36][209], dotarray[37][209], dotarray[38][209], dotarray[39][209], dotarray[40][209], dotarray[41][209], dotarray[42][209], dotarray[43][209], dotarray[44][209], dotarray[45][209], dotarray[46][209], dotarray[47][209], dotarray[48][209], dotarray[49][209], dotarray[50][209], dotarray[51][209], dotarray[52][209], dotarray[53][209], dotarray[54][209], dotarray[55][209], dotarray[56][209], dotarray[57][209], dotarray[58][209], dotarray[59][209], dotarray[60][209], dotarray[61][209], dotarray[62][209], dotarray[63][209], dotarray[64][209], dotarray[65][209], dotarray[66][209], dotarray[67][209], dotarray[68][209], dotarray[69][209], dotarray[70][209], dotarray[71][209], dotarray[72][209], dotarray[73][209], dotarray[74][209], dotarray[75][209], dotarray[76][209], dotarray[77][209], dotarray[78][209], dotarray[79][209], dotarray[80][209], dotarray[81][209], dotarray[82][209], dotarray[83][209], dotarray[84][209], dotarray[85][209], dotarray[86][209], dotarray[87][209], dotarray[88][209], dotarray[89][209], dotarray[90][209], dotarray[91][209], dotarray[92][209], dotarray[93][209], dotarray[94][209], dotarray[95][209], dotarray[96][209], dotarray[97][209], dotarray[98][209], dotarray[99][209], dotarray[100][209], dotarray[101][209], dotarray[102][209], dotarray[103][209], dotarray[104][209], dotarray[105][209], dotarray[106][209], dotarray[107][209], dotarray[108][209], dotarray[109][209], dotarray[110][209], dotarray[111][209], dotarray[112][209], dotarray[113][209], dotarray[114][209], dotarray[115][209], dotarray[116][209], dotarray[117][209], dotarray[118][209], dotarray[119][209], dotarray[120][209], dotarray[121][209], dotarray[122][209], dotarray[123][209], dotarray[124][209], dotarray[125][209], dotarray[126][209], dotarray[127][209]};
assign dot_col_210 = {dotarray[0][210], dotarray[1][210], dotarray[2][210], dotarray[3][210], dotarray[4][210], dotarray[5][210], dotarray[6][210], dotarray[7][210], dotarray[8][210], dotarray[9][210], dotarray[10][210], dotarray[11][210], dotarray[12][210], dotarray[13][210], dotarray[14][210], dotarray[15][210], dotarray[16][210], dotarray[17][210], dotarray[18][210], dotarray[19][210], dotarray[20][210], dotarray[21][210], dotarray[22][210], dotarray[23][210], dotarray[24][210], dotarray[25][210], dotarray[26][210], dotarray[27][210], dotarray[28][210], dotarray[29][210], dotarray[30][210], dotarray[31][210], dotarray[32][210], dotarray[33][210], dotarray[34][210], dotarray[35][210], dotarray[36][210], dotarray[37][210], dotarray[38][210], dotarray[39][210], dotarray[40][210], dotarray[41][210], dotarray[42][210], dotarray[43][210], dotarray[44][210], dotarray[45][210], dotarray[46][210], dotarray[47][210], dotarray[48][210], dotarray[49][210], dotarray[50][210], dotarray[51][210], dotarray[52][210], dotarray[53][210], dotarray[54][210], dotarray[55][210], dotarray[56][210], dotarray[57][210], dotarray[58][210], dotarray[59][210], dotarray[60][210], dotarray[61][210], dotarray[62][210], dotarray[63][210], dotarray[64][210], dotarray[65][210], dotarray[66][210], dotarray[67][210], dotarray[68][210], dotarray[69][210], dotarray[70][210], dotarray[71][210], dotarray[72][210], dotarray[73][210], dotarray[74][210], dotarray[75][210], dotarray[76][210], dotarray[77][210], dotarray[78][210], dotarray[79][210], dotarray[80][210], dotarray[81][210], dotarray[82][210], dotarray[83][210], dotarray[84][210], dotarray[85][210], dotarray[86][210], dotarray[87][210], dotarray[88][210], dotarray[89][210], dotarray[90][210], dotarray[91][210], dotarray[92][210], dotarray[93][210], dotarray[94][210], dotarray[95][210], dotarray[96][210], dotarray[97][210], dotarray[98][210], dotarray[99][210], dotarray[100][210], dotarray[101][210], dotarray[102][210], dotarray[103][210], dotarray[104][210], dotarray[105][210], dotarray[106][210], dotarray[107][210], dotarray[108][210], dotarray[109][210], dotarray[110][210], dotarray[111][210], dotarray[112][210], dotarray[113][210], dotarray[114][210], dotarray[115][210], dotarray[116][210], dotarray[117][210], dotarray[118][210], dotarray[119][210], dotarray[120][210], dotarray[121][210], dotarray[122][210], dotarray[123][210], dotarray[124][210], dotarray[125][210], dotarray[126][210], dotarray[127][210]};
assign dot_col_211 = {dotarray[0][211], dotarray[1][211], dotarray[2][211], dotarray[3][211], dotarray[4][211], dotarray[5][211], dotarray[6][211], dotarray[7][211], dotarray[8][211], dotarray[9][211], dotarray[10][211], dotarray[11][211], dotarray[12][211], dotarray[13][211], dotarray[14][211], dotarray[15][211], dotarray[16][211], dotarray[17][211], dotarray[18][211], dotarray[19][211], dotarray[20][211], dotarray[21][211], dotarray[22][211], dotarray[23][211], dotarray[24][211], dotarray[25][211], dotarray[26][211], dotarray[27][211], dotarray[28][211], dotarray[29][211], dotarray[30][211], dotarray[31][211], dotarray[32][211], dotarray[33][211], dotarray[34][211], dotarray[35][211], dotarray[36][211], dotarray[37][211], dotarray[38][211], dotarray[39][211], dotarray[40][211], dotarray[41][211], dotarray[42][211], dotarray[43][211], dotarray[44][211], dotarray[45][211], dotarray[46][211], dotarray[47][211], dotarray[48][211], dotarray[49][211], dotarray[50][211], dotarray[51][211], dotarray[52][211], dotarray[53][211], dotarray[54][211], dotarray[55][211], dotarray[56][211], dotarray[57][211], dotarray[58][211], dotarray[59][211], dotarray[60][211], dotarray[61][211], dotarray[62][211], dotarray[63][211], dotarray[64][211], dotarray[65][211], dotarray[66][211], dotarray[67][211], dotarray[68][211], dotarray[69][211], dotarray[70][211], dotarray[71][211], dotarray[72][211], dotarray[73][211], dotarray[74][211], dotarray[75][211], dotarray[76][211], dotarray[77][211], dotarray[78][211], dotarray[79][211], dotarray[80][211], dotarray[81][211], dotarray[82][211], dotarray[83][211], dotarray[84][211], dotarray[85][211], dotarray[86][211], dotarray[87][211], dotarray[88][211], dotarray[89][211], dotarray[90][211], dotarray[91][211], dotarray[92][211], dotarray[93][211], dotarray[94][211], dotarray[95][211], dotarray[96][211], dotarray[97][211], dotarray[98][211], dotarray[99][211], dotarray[100][211], dotarray[101][211], dotarray[102][211], dotarray[103][211], dotarray[104][211], dotarray[105][211], dotarray[106][211], dotarray[107][211], dotarray[108][211], dotarray[109][211], dotarray[110][211], dotarray[111][211], dotarray[112][211], dotarray[113][211], dotarray[114][211], dotarray[115][211], dotarray[116][211], dotarray[117][211], dotarray[118][211], dotarray[119][211], dotarray[120][211], dotarray[121][211], dotarray[122][211], dotarray[123][211], dotarray[124][211], dotarray[125][211], dotarray[126][211], dotarray[127][211]};
assign dot_col_212 = {dotarray[0][212], dotarray[1][212], dotarray[2][212], dotarray[3][212], dotarray[4][212], dotarray[5][212], dotarray[6][212], dotarray[7][212], dotarray[8][212], dotarray[9][212], dotarray[10][212], dotarray[11][212], dotarray[12][212], dotarray[13][212], dotarray[14][212], dotarray[15][212], dotarray[16][212], dotarray[17][212], dotarray[18][212], dotarray[19][212], dotarray[20][212], dotarray[21][212], dotarray[22][212], dotarray[23][212], dotarray[24][212], dotarray[25][212], dotarray[26][212], dotarray[27][212], dotarray[28][212], dotarray[29][212], dotarray[30][212], dotarray[31][212], dotarray[32][212], dotarray[33][212], dotarray[34][212], dotarray[35][212], dotarray[36][212], dotarray[37][212], dotarray[38][212], dotarray[39][212], dotarray[40][212], dotarray[41][212], dotarray[42][212], dotarray[43][212], dotarray[44][212], dotarray[45][212], dotarray[46][212], dotarray[47][212], dotarray[48][212], dotarray[49][212], dotarray[50][212], dotarray[51][212], dotarray[52][212], dotarray[53][212], dotarray[54][212], dotarray[55][212], dotarray[56][212], dotarray[57][212], dotarray[58][212], dotarray[59][212], dotarray[60][212], dotarray[61][212], dotarray[62][212], dotarray[63][212], dotarray[64][212], dotarray[65][212], dotarray[66][212], dotarray[67][212], dotarray[68][212], dotarray[69][212], dotarray[70][212], dotarray[71][212], dotarray[72][212], dotarray[73][212], dotarray[74][212], dotarray[75][212], dotarray[76][212], dotarray[77][212], dotarray[78][212], dotarray[79][212], dotarray[80][212], dotarray[81][212], dotarray[82][212], dotarray[83][212], dotarray[84][212], dotarray[85][212], dotarray[86][212], dotarray[87][212], dotarray[88][212], dotarray[89][212], dotarray[90][212], dotarray[91][212], dotarray[92][212], dotarray[93][212], dotarray[94][212], dotarray[95][212], dotarray[96][212], dotarray[97][212], dotarray[98][212], dotarray[99][212], dotarray[100][212], dotarray[101][212], dotarray[102][212], dotarray[103][212], dotarray[104][212], dotarray[105][212], dotarray[106][212], dotarray[107][212], dotarray[108][212], dotarray[109][212], dotarray[110][212], dotarray[111][212], dotarray[112][212], dotarray[113][212], dotarray[114][212], dotarray[115][212], dotarray[116][212], dotarray[117][212], dotarray[118][212], dotarray[119][212], dotarray[120][212], dotarray[121][212], dotarray[122][212], dotarray[123][212], dotarray[124][212], dotarray[125][212], dotarray[126][212], dotarray[127][212]};
assign dot_col_213 = {dotarray[0][213], dotarray[1][213], dotarray[2][213], dotarray[3][213], dotarray[4][213], dotarray[5][213], dotarray[6][213], dotarray[7][213], dotarray[8][213], dotarray[9][213], dotarray[10][213], dotarray[11][213], dotarray[12][213], dotarray[13][213], dotarray[14][213], dotarray[15][213], dotarray[16][213], dotarray[17][213], dotarray[18][213], dotarray[19][213], dotarray[20][213], dotarray[21][213], dotarray[22][213], dotarray[23][213], dotarray[24][213], dotarray[25][213], dotarray[26][213], dotarray[27][213], dotarray[28][213], dotarray[29][213], dotarray[30][213], dotarray[31][213], dotarray[32][213], dotarray[33][213], dotarray[34][213], dotarray[35][213], dotarray[36][213], dotarray[37][213], dotarray[38][213], dotarray[39][213], dotarray[40][213], dotarray[41][213], dotarray[42][213], dotarray[43][213], dotarray[44][213], dotarray[45][213], dotarray[46][213], dotarray[47][213], dotarray[48][213], dotarray[49][213], dotarray[50][213], dotarray[51][213], dotarray[52][213], dotarray[53][213], dotarray[54][213], dotarray[55][213], dotarray[56][213], dotarray[57][213], dotarray[58][213], dotarray[59][213], dotarray[60][213], dotarray[61][213], dotarray[62][213], dotarray[63][213], dotarray[64][213], dotarray[65][213], dotarray[66][213], dotarray[67][213], dotarray[68][213], dotarray[69][213], dotarray[70][213], dotarray[71][213], dotarray[72][213], dotarray[73][213], dotarray[74][213], dotarray[75][213], dotarray[76][213], dotarray[77][213], dotarray[78][213], dotarray[79][213], dotarray[80][213], dotarray[81][213], dotarray[82][213], dotarray[83][213], dotarray[84][213], dotarray[85][213], dotarray[86][213], dotarray[87][213], dotarray[88][213], dotarray[89][213], dotarray[90][213], dotarray[91][213], dotarray[92][213], dotarray[93][213], dotarray[94][213], dotarray[95][213], dotarray[96][213], dotarray[97][213], dotarray[98][213], dotarray[99][213], dotarray[100][213], dotarray[101][213], dotarray[102][213], dotarray[103][213], dotarray[104][213], dotarray[105][213], dotarray[106][213], dotarray[107][213], dotarray[108][213], dotarray[109][213], dotarray[110][213], dotarray[111][213], dotarray[112][213], dotarray[113][213], dotarray[114][213], dotarray[115][213], dotarray[116][213], dotarray[117][213], dotarray[118][213], dotarray[119][213], dotarray[120][213], dotarray[121][213], dotarray[122][213], dotarray[123][213], dotarray[124][213], dotarray[125][213], dotarray[126][213], dotarray[127][213]};
assign dot_col_214 = {dotarray[0][214], dotarray[1][214], dotarray[2][214], dotarray[3][214], dotarray[4][214], dotarray[5][214], dotarray[6][214], dotarray[7][214], dotarray[8][214], dotarray[9][214], dotarray[10][214], dotarray[11][214], dotarray[12][214], dotarray[13][214], dotarray[14][214], dotarray[15][214], dotarray[16][214], dotarray[17][214], dotarray[18][214], dotarray[19][214], dotarray[20][214], dotarray[21][214], dotarray[22][214], dotarray[23][214], dotarray[24][214], dotarray[25][214], dotarray[26][214], dotarray[27][214], dotarray[28][214], dotarray[29][214], dotarray[30][214], dotarray[31][214], dotarray[32][214], dotarray[33][214], dotarray[34][214], dotarray[35][214], dotarray[36][214], dotarray[37][214], dotarray[38][214], dotarray[39][214], dotarray[40][214], dotarray[41][214], dotarray[42][214], dotarray[43][214], dotarray[44][214], dotarray[45][214], dotarray[46][214], dotarray[47][214], dotarray[48][214], dotarray[49][214], dotarray[50][214], dotarray[51][214], dotarray[52][214], dotarray[53][214], dotarray[54][214], dotarray[55][214], dotarray[56][214], dotarray[57][214], dotarray[58][214], dotarray[59][214], dotarray[60][214], dotarray[61][214], dotarray[62][214], dotarray[63][214], dotarray[64][214], dotarray[65][214], dotarray[66][214], dotarray[67][214], dotarray[68][214], dotarray[69][214], dotarray[70][214], dotarray[71][214], dotarray[72][214], dotarray[73][214], dotarray[74][214], dotarray[75][214], dotarray[76][214], dotarray[77][214], dotarray[78][214], dotarray[79][214], dotarray[80][214], dotarray[81][214], dotarray[82][214], dotarray[83][214], dotarray[84][214], dotarray[85][214], dotarray[86][214], dotarray[87][214], dotarray[88][214], dotarray[89][214], dotarray[90][214], dotarray[91][214], dotarray[92][214], dotarray[93][214], dotarray[94][214], dotarray[95][214], dotarray[96][214], dotarray[97][214], dotarray[98][214], dotarray[99][214], dotarray[100][214], dotarray[101][214], dotarray[102][214], dotarray[103][214], dotarray[104][214], dotarray[105][214], dotarray[106][214], dotarray[107][214], dotarray[108][214], dotarray[109][214], dotarray[110][214], dotarray[111][214], dotarray[112][214], dotarray[113][214], dotarray[114][214], dotarray[115][214], dotarray[116][214], dotarray[117][214], dotarray[118][214], dotarray[119][214], dotarray[120][214], dotarray[121][214], dotarray[122][214], dotarray[123][214], dotarray[124][214], dotarray[125][214], dotarray[126][214], dotarray[127][214]};
assign dot_col_215 = {dotarray[0][215], dotarray[1][215], dotarray[2][215], dotarray[3][215], dotarray[4][215], dotarray[5][215], dotarray[6][215], dotarray[7][215], dotarray[8][215], dotarray[9][215], dotarray[10][215], dotarray[11][215], dotarray[12][215], dotarray[13][215], dotarray[14][215], dotarray[15][215], dotarray[16][215], dotarray[17][215], dotarray[18][215], dotarray[19][215], dotarray[20][215], dotarray[21][215], dotarray[22][215], dotarray[23][215], dotarray[24][215], dotarray[25][215], dotarray[26][215], dotarray[27][215], dotarray[28][215], dotarray[29][215], dotarray[30][215], dotarray[31][215], dotarray[32][215], dotarray[33][215], dotarray[34][215], dotarray[35][215], dotarray[36][215], dotarray[37][215], dotarray[38][215], dotarray[39][215], dotarray[40][215], dotarray[41][215], dotarray[42][215], dotarray[43][215], dotarray[44][215], dotarray[45][215], dotarray[46][215], dotarray[47][215], dotarray[48][215], dotarray[49][215], dotarray[50][215], dotarray[51][215], dotarray[52][215], dotarray[53][215], dotarray[54][215], dotarray[55][215], dotarray[56][215], dotarray[57][215], dotarray[58][215], dotarray[59][215], dotarray[60][215], dotarray[61][215], dotarray[62][215], dotarray[63][215], dotarray[64][215], dotarray[65][215], dotarray[66][215], dotarray[67][215], dotarray[68][215], dotarray[69][215], dotarray[70][215], dotarray[71][215], dotarray[72][215], dotarray[73][215], dotarray[74][215], dotarray[75][215], dotarray[76][215], dotarray[77][215], dotarray[78][215], dotarray[79][215], dotarray[80][215], dotarray[81][215], dotarray[82][215], dotarray[83][215], dotarray[84][215], dotarray[85][215], dotarray[86][215], dotarray[87][215], dotarray[88][215], dotarray[89][215], dotarray[90][215], dotarray[91][215], dotarray[92][215], dotarray[93][215], dotarray[94][215], dotarray[95][215], dotarray[96][215], dotarray[97][215], dotarray[98][215], dotarray[99][215], dotarray[100][215], dotarray[101][215], dotarray[102][215], dotarray[103][215], dotarray[104][215], dotarray[105][215], dotarray[106][215], dotarray[107][215], dotarray[108][215], dotarray[109][215], dotarray[110][215], dotarray[111][215], dotarray[112][215], dotarray[113][215], dotarray[114][215], dotarray[115][215], dotarray[116][215], dotarray[117][215], dotarray[118][215], dotarray[119][215], dotarray[120][215], dotarray[121][215], dotarray[122][215], dotarray[123][215], dotarray[124][215], dotarray[125][215], dotarray[126][215], dotarray[127][215]};
assign dot_col_216 = {dotarray[0][216], dotarray[1][216], dotarray[2][216], dotarray[3][216], dotarray[4][216], dotarray[5][216], dotarray[6][216], dotarray[7][216], dotarray[8][216], dotarray[9][216], dotarray[10][216], dotarray[11][216], dotarray[12][216], dotarray[13][216], dotarray[14][216], dotarray[15][216], dotarray[16][216], dotarray[17][216], dotarray[18][216], dotarray[19][216], dotarray[20][216], dotarray[21][216], dotarray[22][216], dotarray[23][216], dotarray[24][216], dotarray[25][216], dotarray[26][216], dotarray[27][216], dotarray[28][216], dotarray[29][216], dotarray[30][216], dotarray[31][216], dotarray[32][216], dotarray[33][216], dotarray[34][216], dotarray[35][216], dotarray[36][216], dotarray[37][216], dotarray[38][216], dotarray[39][216], dotarray[40][216], dotarray[41][216], dotarray[42][216], dotarray[43][216], dotarray[44][216], dotarray[45][216], dotarray[46][216], dotarray[47][216], dotarray[48][216], dotarray[49][216], dotarray[50][216], dotarray[51][216], dotarray[52][216], dotarray[53][216], dotarray[54][216], dotarray[55][216], dotarray[56][216], dotarray[57][216], dotarray[58][216], dotarray[59][216], dotarray[60][216], dotarray[61][216], dotarray[62][216], dotarray[63][216], dotarray[64][216], dotarray[65][216], dotarray[66][216], dotarray[67][216], dotarray[68][216], dotarray[69][216], dotarray[70][216], dotarray[71][216], dotarray[72][216], dotarray[73][216], dotarray[74][216], dotarray[75][216], dotarray[76][216], dotarray[77][216], dotarray[78][216], dotarray[79][216], dotarray[80][216], dotarray[81][216], dotarray[82][216], dotarray[83][216], dotarray[84][216], dotarray[85][216], dotarray[86][216], dotarray[87][216], dotarray[88][216], dotarray[89][216], dotarray[90][216], dotarray[91][216], dotarray[92][216], dotarray[93][216], dotarray[94][216], dotarray[95][216], dotarray[96][216], dotarray[97][216], dotarray[98][216], dotarray[99][216], dotarray[100][216], dotarray[101][216], dotarray[102][216], dotarray[103][216], dotarray[104][216], dotarray[105][216], dotarray[106][216], dotarray[107][216], dotarray[108][216], dotarray[109][216], dotarray[110][216], dotarray[111][216], dotarray[112][216], dotarray[113][216], dotarray[114][216], dotarray[115][216], dotarray[116][216], dotarray[117][216], dotarray[118][216], dotarray[119][216], dotarray[120][216], dotarray[121][216], dotarray[122][216], dotarray[123][216], dotarray[124][216], dotarray[125][216], dotarray[126][216], dotarray[127][216]};
assign dot_col_217 = {dotarray[0][217], dotarray[1][217], dotarray[2][217], dotarray[3][217], dotarray[4][217], dotarray[5][217], dotarray[6][217], dotarray[7][217], dotarray[8][217], dotarray[9][217], dotarray[10][217], dotarray[11][217], dotarray[12][217], dotarray[13][217], dotarray[14][217], dotarray[15][217], dotarray[16][217], dotarray[17][217], dotarray[18][217], dotarray[19][217], dotarray[20][217], dotarray[21][217], dotarray[22][217], dotarray[23][217], dotarray[24][217], dotarray[25][217], dotarray[26][217], dotarray[27][217], dotarray[28][217], dotarray[29][217], dotarray[30][217], dotarray[31][217], dotarray[32][217], dotarray[33][217], dotarray[34][217], dotarray[35][217], dotarray[36][217], dotarray[37][217], dotarray[38][217], dotarray[39][217], dotarray[40][217], dotarray[41][217], dotarray[42][217], dotarray[43][217], dotarray[44][217], dotarray[45][217], dotarray[46][217], dotarray[47][217], dotarray[48][217], dotarray[49][217], dotarray[50][217], dotarray[51][217], dotarray[52][217], dotarray[53][217], dotarray[54][217], dotarray[55][217], dotarray[56][217], dotarray[57][217], dotarray[58][217], dotarray[59][217], dotarray[60][217], dotarray[61][217], dotarray[62][217], dotarray[63][217], dotarray[64][217], dotarray[65][217], dotarray[66][217], dotarray[67][217], dotarray[68][217], dotarray[69][217], dotarray[70][217], dotarray[71][217], dotarray[72][217], dotarray[73][217], dotarray[74][217], dotarray[75][217], dotarray[76][217], dotarray[77][217], dotarray[78][217], dotarray[79][217], dotarray[80][217], dotarray[81][217], dotarray[82][217], dotarray[83][217], dotarray[84][217], dotarray[85][217], dotarray[86][217], dotarray[87][217], dotarray[88][217], dotarray[89][217], dotarray[90][217], dotarray[91][217], dotarray[92][217], dotarray[93][217], dotarray[94][217], dotarray[95][217], dotarray[96][217], dotarray[97][217], dotarray[98][217], dotarray[99][217], dotarray[100][217], dotarray[101][217], dotarray[102][217], dotarray[103][217], dotarray[104][217], dotarray[105][217], dotarray[106][217], dotarray[107][217], dotarray[108][217], dotarray[109][217], dotarray[110][217], dotarray[111][217], dotarray[112][217], dotarray[113][217], dotarray[114][217], dotarray[115][217], dotarray[116][217], dotarray[117][217], dotarray[118][217], dotarray[119][217], dotarray[120][217], dotarray[121][217], dotarray[122][217], dotarray[123][217], dotarray[124][217], dotarray[125][217], dotarray[126][217], dotarray[127][217]};
assign dot_col_218 = {dotarray[0][218], dotarray[1][218], dotarray[2][218], dotarray[3][218], dotarray[4][218], dotarray[5][218], dotarray[6][218], dotarray[7][218], dotarray[8][218], dotarray[9][218], dotarray[10][218], dotarray[11][218], dotarray[12][218], dotarray[13][218], dotarray[14][218], dotarray[15][218], dotarray[16][218], dotarray[17][218], dotarray[18][218], dotarray[19][218], dotarray[20][218], dotarray[21][218], dotarray[22][218], dotarray[23][218], dotarray[24][218], dotarray[25][218], dotarray[26][218], dotarray[27][218], dotarray[28][218], dotarray[29][218], dotarray[30][218], dotarray[31][218], dotarray[32][218], dotarray[33][218], dotarray[34][218], dotarray[35][218], dotarray[36][218], dotarray[37][218], dotarray[38][218], dotarray[39][218], dotarray[40][218], dotarray[41][218], dotarray[42][218], dotarray[43][218], dotarray[44][218], dotarray[45][218], dotarray[46][218], dotarray[47][218], dotarray[48][218], dotarray[49][218], dotarray[50][218], dotarray[51][218], dotarray[52][218], dotarray[53][218], dotarray[54][218], dotarray[55][218], dotarray[56][218], dotarray[57][218], dotarray[58][218], dotarray[59][218], dotarray[60][218], dotarray[61][218], dotarray[62][218], dotarray[63][218], dotarray[64][218], dotarray[65][218], dotarray[66][218], dotarray[67][218], dotarray[68][218], dotarray[69][218], dotarray[70][218], dotarray[71][218], dotarray[72][218], dotarray[73][218], dotarray[74][218], dotarray[75][218], dotarray[76][218], dotarray[77][218], dotarray[78][218], dotarray[79][218], dotarray[80][218], dotarray[81][218], dotarray[82][218], dotarray[83][218], dotarray[84][218], dotarray[85][218], dotarray[86][218], dotarray[87][218], dotarray[88][218], dotarray[89][218], dotarray[90][218], dotarray[91][218], dotarray[92][218], dotarray[93][218], dotarray[94][218], dotarray[95][218], dotarray[96][218], dotarray[97][218], dotarray[98][218], dotarray[99][218], dotarray[100][218], dotarray[101][218], dotarray[102][218], dotarray[103][218], dotarray[104][218], dotarray[105][218], dotarray[106][218], dotarray[107][218], dotarray[108][218], dotarray[109][218], dotarray[110][218], dotarray[111][218], dotarray[112][218], dotarray[113][218], dotarray[114][218], dotarray[115][218], dotarray[116][218], dotarray[117][218], dotarray[118][218], dotarray[119][218], dotarray[120][218], dotarray[121][218], dotarray[122][218], dotarray[123][218], dotarray[124][218], dotarray[125][218], dotarray[126][218], dotarray[127][218]};
assign dot_col_219 = {dotarray[0][219], dotarray[1][219], dotarray[2][219], dotarray[3][219], dotarray[4][219], dotarray[5][219], dotarray[6][219], dotarray[7][219], dotarray[8][219], dotarray[9][219], dotarray[10][219], dotarray[11][219], dotarray[12][219], dotarray[13][219], dotarray[14][219], dotarray[15][219], dotarray[16][219], dotarray[17][219], dotarray[18][219], dotarray[19][219], dotarray[20][219], dotarray[21][219], dotarray[22][219], dotarray[23][219], dotarray[24][219], dotarray[25][219], dotarray[26][219], dotarray[27][219], dotarray[28][219], dotarray[29][219], dotarray[30][219], dotarray[31][219], dotarray[32][219], dotarray[33][219], dotarray[34][219], dotarray[35][219], dotarray[36][219], dotarray[37][219], dotarray[38][219], dotarray[39][219], dotarray[40][219], dotarray[41][219], dotarray[42][219], dotarray[43][219], dotarray[44][219], dotarray[45][219], dotarray[46][219], dotarray[47][219], dotarray[48][219], dotarray[49][219], dotarray[50][219], dotarray[51][219], dotarray[52][219], dotarray[53][219], dotarray[54][219], dotarray[55][219], dotarray[56][219], dotarray[57][219], dotarray[58][219], dotarray[59][219], dotarray[60][219], dotarray[61][219], dotarray[62][219], dotarray[63][219], dotarray[64][219], dotarray[65][219], dotarray[66][219], dotarray[67][219], dotarray[68][219], dotarray[69][219], dotarray[70][219], dotarray[71][219], dotarray[72][219], dotarray[73][219], dotarray[74][219], dotarray[75][219], dotarray[76][219], dotarray[77][219], dotarray[78][219], dotarray[79][219], dotarray[80][219], dotarray[81][219], dotarray[82][219], dotarray[83][219], dotarray[84][219], dotarray[85][219], dotarray[86][219], dotarray[87][219], dotarray[88][219], dotarray[89][219], dotarray[90][219], dotarray[91][219], dotarray[92][219], dotarray[93][219], dotarray[94][219], dotarray[95][219], dotarray[96][219], dotarray[97][219], dotarray[98][219], dotarray[99][219], dotarray[100][219], dotarray[101][219], dotarray[102][219], dotarray[103][219], dotarray[104][219], dotarray[105][219], dotarray[106][219], dotarray[107][219], dotarray[108][219], dotarray[109][219], dotarray[110][219], dotarray[111][219], dotarray[112][219], dotarray[113][219], dotarray[114][219], dotarray[115][219], dotarray[116][219], dotarray[117][219], dotarray[118][219], dotarray[119][219], dotarray[120][219], dotarray[121][219], dotarray[122][219], dotarray[123][219], dotarray[124][219], dotarray[125][219], dotarray[126][219], dotarray[127][219]};
assign dot_col_220 = {dotarray[0][220], dotarray[1][220], dotarray[2][220], dotarray[3][220], dotarray[4][220], dotarray[5][220], dotarray[6][220], dotarray[7][220], dotarray[8][220], dotarray[9][220], dotarray[10][220], dotarray[11][220], dotarray[12][220], dotarray[13][220], dotarray[14][220], dotarray[15][220], dotarray[16][220], dotarray[17][220], dotarray[18][220], dotarray[19][220], dotarray[20][220], dotarray[21][220], dotarray[22][220], dotarray[23][220], dotarray[24][220], dotarray[25][220], dotarray[26][220], dotarray[27][220], dotarray[28][220], dotarray[29][220], dotarray[30][220], dotarray[31][220], dotarray[32][220], dotarray[33][220], dotarray[34][220], dotarray[35][220], dotarray[36][220], dotarray[37][220], dotarray[38][220], dotarray[39][220], dotarray[40][220], dotarray[41][220], dotarray[42][220], dotarray[43][220], dotarray[44][220], dotarray[45][220], dotarray[46][220], dotarray[47][220], dotarray[48][220], dotarray[49][220], dotarray[50][220], dotarray[51][220], dotarray[52][220], dotarray[53][220], dotarray[54][220], dotarray[55][220], dotarray[56][220], dotarray[57][220], dotarray[58][220], dotarray[59][220], dotarray[60][220], dotarray[61][220], dotarray[62][220], dotarray[63][220], dotarray[64][220], dotarray[65][220], dotarray[66][220], dotarray[67][220], dotarray[68][220], dotarray[69][220], dotarray[70][220], dotarray[71][220], dotarray[72][220], dotarray[73][220], dotarray[74][220], dotarray[75][220], dotarray[76][220], dotarray[77][220], dotarray[78][220], dotarray[79][220], dotarray[80][220], dotarray[81][220], dotarray[82][220], dotarray[83][220], dotarray[84][220], dotarray[85][220], dotarray[86][220], dotarray[87][220], dotarray[88][220], dotarray[89][220], dotarray[90][220], dotarray[91][220], dotarray[92][220], dotarray[93][220], dotarray[94][220], dotarray[95][220], dotarray[96][220], dotarray[97][220], dotarray[98][220], dotarray[99][220], dotarray[100][220], dotarray[101][220], dotarray[102][220], dotarray[103][220], dotarray[104][220], dotarray[105][220], dotarray[106][220], dotarray[107][220], dotarray[108][220], dotarray[109][220], dotarray[110][220], dotarray[111][220], dotarray[112][220], dotarray[113][220], dotarray[114][220], dotarray[115][220], dotarray[116][220], dotarray[117][220], dotarray[118][220], dotarray[119][220], dotarray[120][220], dotarray[121][220], dotarray[122][220], dotarray[123][220], dotarray[124][220], dotarray[125][220], dotarray[126][220], dotarray[127][220]};
assign dot_col_221 = {dotarray[0][221], dotarray[1][221], dotarray[2][221], dotarray[3][221], dotarray[4][221], dotarray[5][221], dotarray[6][221], dotarray[7][221], dotarray[8][221], dotarray[9][221], dotarray[10][221], dotarray[11][221], dotarray[12][221], dotarray[13][221], dotarray[14][221], dotarray[15][221], dotarray[16][221], dotarray[17][221], dotarray[18][221], dotarray[19][221], dotarray[20][221], dotarray[21][221], dotarray[22][221], dotarray[23][221], dotarray[24][221], dotarray[25][221], dotarray[26][221], dotarray[27][221], dotarray[28][221], dotarray[29][221], dotarray[30][221], dotarray[31][221], dotarray[32][221], dotarray[33][221], dotarray[34][221], dotarray[35][221], dotarray[36][221], dotarray[37][221], dotarray[38][221], dotarray[39][221], dotarray[40][221], dotarray[41][221], dotarray[42][221], dotarray[43][221], dotarray[44][221], dotarray[45][221], dotarray[46][221], dotarray[47][221], dotarray[48][221], dotarray[49][221], dotarray[50][221], dotarray[51][221], dotarray[52][221], dotarray[53][221], dotarray[54][221], dotarray[55][221], dotarray[56][221], dotarray[57][221], dotarray[58][221], dotarray[59][221], dotarray[60][221], dotarray[61][221], dotarray[62][221], dotarray[63][221], dotarray[64][221], dotarray[65][221], dotarray[66][221], dotarray[67][221], dotarray[68][221], dotarray[69][221], dotarray[70][221], dotarray[71][221], dotarray[72][221], dotarray[73][221], dotarray[74][221], dotarray[75][221], dotarray[76][221], dotarray[77][221], dotarray[78][221], dotarray[79][221], dotarray[80][221], dotarray[81][221], dotarray[82][221], dotarray[83][221], dotarray[84][221], dotarray[85][221], dotarray[86][221], dotarray[87][221], dotarray[88][221], dotarray[89][221], dotarray[90][221], dotarray[91][221], dotarray[92][221], dotarray[93][221], dotarray[94][221], dotarray[95][221], dotarray[96][221], dotarray[97][221], dotarray[98][221], dotarray[99][221], dotarray[100][221], dotarray[101][221], dotarray[102][221], dotarray[103][221], dotarray[104][221], dotarray[105][221], dotarray[106][221], dotarray[107][221], dotarray[108][221], dotarray[109][221], dotarray[110][221], dotarray[111][221], dotarray[112][221], dotarray[113][221], dotarray[114][221], dotarray[115][221], dotarray[116][221], dotarray[117][221], dotarray[118][221], dotarray[119][221], dotarray[120][221], dotarray[121][221], dotarray[122][221], dotarray[123][221], dotarray[124][221], dotarray[125][221], dotarray[126][221], dotarray[127][221]};
assign dot_col_222 = {dotarray[0][222], dotarray[1][222], dotarray[2][222], dotarray[3][222], dotarray[4][222], dotarray[5][222], dotarray[6][222], dotarray[7][222], dotarray[8][222], dotarray[9][222], dotarray[10][222], dotarray[11][222], dotarray[12][222], dotarray[13][222], dotarray[14][222], dotarray[15][222], dotarray[16][222], dotarray[17][222], dotarray[18][222], dotarray[19][222], dotarray[20][222], dotarray[21][222], dotarray[22][222], dotarray[23][222], dotarray[24][222], dotarray[25][222], dotarray[26][222], dotarray[27][222], dotarray[28][222], dotarray[29][222], dotarray[30][222], dotarray[31][222], dotarray[32][222], dotarray[33][222], dotarray[34][222], dotarray[35][222], dotarray[36][222], dotarray[37][222], dotarray[38][222], dotarray[39][222], dotarray[40][222], dotarray[41][222], dotarray[42][222], dotarray[43][222], dotarray[44][222], dotarray[45][222], dotarray[46][222], dotarray[47][222], dotarray[48][222], dotarray[49][222], dotarray[50][222], dotarray[51][222], dotarray[52][222], dotarray[53][222], dotarray[54][222], dotarray[55][222], dotarray[56][222], dotarray[57][222], dotarray[58][222], dotarray[59][222], dotarray[60][222], dotarray[61][222], dotarray[62][222], dotarray[63][222], dotarray[64][222], dotarray[65][222], dotarray[66][222], dotarray[67][222], dotarray[68][222], dotarray[69][222], dotarray[70][222], dotarray[71][222], dotarray[72][222], dotarray[73][222], dotarray[74][222], dotarray[75][222], dotarray[76][222], dotarray[77][222], dotarray[78][222], dotarray[79][222], dotarray[80][222], dotarray[81][222], dotarray[82][222], dotarray[83][222], dotarray[84][222], dotarray[85][222], dotarray[86][222], dotarray[87][222], dotarray[88][222], dotarray[89][222], dotarray[90][222], dotarray[91][222], dotarray[92][222], dotarray[93][222], dotarray[94][222], dotarray[95][222], dotarray[96][222], dotarray[97][222], dotarray[98][222], dotarray[99][222], dotarray[100][222], dotarray[101][222], dotarray[102][222], dotarray[103][222], dotarray[104][222], dotarray[105][222], dotarray[106][222], dotarray[107][222], dotarray[108][222], dotarray[109][222], dotarray[110][222], dotarray[111][222], dotarray[112][222], dotarray[113][222], dotarray[114][222], dotarray[115][222], dotarray[116][222], dotarray[117][222], dotarray[118][222], dotarray[119][222], dotarray[120][222], dotarray[121][222], dotarray[122][222], dotarray[123][222], dotarray[124][222], dotarray[125][222], dotarray[126][222], dotarray[127][222]};
assign dot_col_223 = {dotarray[0][223], dotarray[1][223], dotarray[2][223], dotarray[3][223], dotarray[4][223], dotarray[5][223], dotarray[6][223], dotarray[7][223], dotarray[8][223], dotarray[9][223], dotarray[10][223], dotarray[11][223], dotarray[12][223], dotarray[13][223], dotarray[14][223], dotarray[15][223], dotarray[16][223], dotarray[17][223], dotarray[18][223], dotarray[19][223], dotarray[20][223], dotarray[21][223], dotarray[22][223], dotarray[23][223], dotarray[24][223], dotarray[25][223], dotarray[26][223], dotarray[27][223], dotarray[28][223], dotarray[29][223], dotarray[30][223], dotarray[31][223], dotarray[32][223], dotarray[33][223], dotarray[34][223], dotarray[35][223], dotarray[36][223], dotarray[37][223], dotarray[38][223], dotarray[39][223], dotarray[40][223], dotarray[41][223], dotarray[42][223], dotarray[43][223], dotarray[44][223], dotarray[45][223], dotarray[46][223], dotarray[47][223], dotarray[48][223], dotarray[49][223], dotarray[50][223], dotarray[51][223], dotarray[52][223], dotarray[53][223], dotarray[54][223], dotarray[55][223], dotarray[56][223], dotarray[57][223], dotarray[58][223], dotarray[59][223], dotarray[60][223], dotarray[61][223], dotarray[62][223], dotarray[63][223], dotarray[64][223], dotarray[65][223], dotarray[66][223], dotarray[67][223], dotarray[68][223], dotarray[69][223], dotarray[70][223], dotarray[71][223], dotarray[72][223], dotarray[73][223], dotarray[74][223], dotarray[75][223], dotarray[76][223], dotarray[77][223], dotarray[78][223], dotarray[79][223], dotarray[80][223], dotarray[81][223], dotarray[82][223], dotarray[83][223], dotarray[84][223], dotarray[85][223], dotarray[86][223], dotarray[87][223], dotarray[88][223], dotarray[89][223], dotarray[90][223], dotarray[91][223], dotarray[92][223], dotarray[93][223], dotarray[94][223], dotarray[95][223], dotarray[96][223], dotarray[97][223], dotarray[98][223], dotarray[99][223], dotarray[100][223], dotarray[101][223], dotarray[102][223], dotarray[103][223], dotarray[104][223], dotarray[105][223], dotarray[106][223], dotarray[107][223], dotarray[108][223], dotarray[109][223], dotarray[110][223], dotarray[111][223], dotarray[112][223], dotarray[113][223], dotarray[114][223], dotarray[115][223], dotarray[116][223], dotarray[117][223], dotarray[118][223], dotarray[119][223], dotarray[120][223], dotarray[121][223], dotarray[122][223], dotarray[123][223], dotarray[124][223], dotarray[125][223], dotarray[126][223], dotarray[127][223]};
assign dot_col_224 = {dotarray[0][224], dotarray[1][224], dotarray[2][224], dotarray[3][224], dotarray[4][224], dotarray[5][224], dotarray[6][224], dotarray[7][224], dotarray[8][224], dotarray[9][224], dotarray[10][224], dotarray[11][224], dotarray[12][224], dotarray[13][224], dotarray[14][224], dotarray[15][224], dotarray[16][224], dotarray[17][224], dotarray[18][224], dotarray[19][224], dotarray[20][224], dotarray[21][224], dotarray[22][224], dotarray[23][224], dotarray[24][224], dotarray[25][224], dotarray[26][224], dotarray[27][224], dotarray[28][224], dotarray[29][224], dotarray[30][224], dotarray[31][224], dotarray[32][224], dotarray[33][224], dotarray[34][224], dotarray[35][224], dotarray[36][224], dotarray[37][224], dotarray[38][224], dotarray[39][224], dotarray[40][224], dotarray[41][224], dotarray[42][224], dotarray[43][224], dotarray[44][224], dotarray[45][224], dotarray[46][224], dotarray[47][224], dotarray[48][224], dotarray[49][224], dotarray[50][224], dotarray[51][224], dotarray[52][224], dotarray[53][224], dotarray[54][224], dotarray[55][224], dotarray[56][224], dotarray[57][224], dotarray[58][224], dotarray[59][224], dotarray[60][224], dotarray[61][224], dotarray[62][224], dotarray[63][224], dotarray[64][224], dotarray[65][224], dotarray[66][224], dotarray[67][224], dotarray[68][224], dotarray[69][224], dotarray[70][224], dotarray[71][224], dotarray[72][224], dotarray[73][224], dotarray[74][224], dotarray[75][224], dotarray[76][224], dotarray[77][224], dotarray[78][224], dotarray[79][224], dotarray[80][224], dotarray[81][224], dotarray[82][224], dotarray[83][224], dotarray[84][224], dotarray[85][224], dotarray[86][224], dotarray[87][224], dotarray[88][224], dotarray[89][224], dotarray[90][224], dotarray[91][224], dotarray[92][224], dotarray[93][224], dotarray[94][224], dotarray[95][224], dotarray[96][224], dotarray[97][224], dotarray[98][224], dotarray[99][224], dotarray[100][224], dotarray[101][224], dotarray[102][224], dotarray[103][224], dotarray[104][224], dotarray[105][224], dotarray[106][224], dotarray[107][224], dotarray[108][224], dotarray[109][224], dotarray[110][224], dotarray[111][224], dotarray[112][224], dotarray[113][224], dotarray[114][224], dotarray[115][224], dotarray[116][224], dotarray[117][224], dotarray[118][224], dotarray[119][224], dotarray[120][224], dotarray[121][224], dotarray[122][224], dotarray[123][224], dotarray[124][224], dotarray[125][224], dotarray[126][224], dotarray[127][224]};
assign dot_col_225 = {dotarray[0][225], dotarray[1][225], dotarray[2][225], dotarray[3][225], dotarray[4][225], dotarray[5][225], dotarray[6][225], dotarray[7][225], dotarray[8][225], dotarray[9][225], dotarray[10][225], dotarray[11][225], dotarray[12][225], dotarray[13][225], dotarray[14][225], dotarray[15][225], dotarray[16][225], dotarray[17][225], dotarray[18][225], dotarray[19][225], dotarray[20][225], dotarray[21][225], dotarray[22][225], dotarray[23][225], dotarray[24][225], dotarray[25][225], dotarray[26][225], dotarray[27][225], dotarray[28][225], dotarray[29][225], dotarray[30][225], dotarray[31][225], dotarray[32][225], dotarray[33][225], dotarray[34][225], dotarray[35][225], dotarray[36][225], dotarray[37][225], dotarray[38][225], dotarray[39][225], dotarray[40][225], dotarray[41][225], dotarray[42][225], dotarray[43][225], dotarray[44][225], dotarray[45][225], dotarray[46][225], dotarray[47][225], dotarray[48][225], dotarray[49][225], dotarray[50][225], dotarray[51][225], dotarray[52][225], dotarray[53][225], dotarray[54][225], dotarray[55][225], dotarray[56][225], dotarray[57][225], dotarray[58][225], dotarray[59][225], dotarray[60][225], dotarray[61][225], dotarray[62][225], dotarray[63][225], dotarray[64][225], dotarray[65][225], dotarray[66][225], dotarray[67][225], dotarray[68][225], dotarray[69][225], dotarray[70][225], dotarray[71][225], dotarray[72][225], dotarray[73][225], dotarray[74][225], dotarray[75][225], dotarray[76][225], dotarray[77][225], dotarray[78][225], dotarray[79][225], dotarray[80][225], dotarray[81][225], dotarray[82][225], dotarray[83][225], dotarray[84][225], dotarray[85][225], dotarray[86][225], dotarray[87][225], dotarray[88][225], dotarray[89][225], dotarray[90][225], dotarray[91][225], dotarray[92][225], dotarray[93][225], dotarray[94][225], dotarray[95][225], dotarray[96][225], dotarray[97][225], dotarray[98][225], dotarray[99][225], dotarray[100][225], dotarray[101][225], dotarray[102][225], dotarray[103][225], dotarray[104][225], dotarray[105][225], dotarray[106][225], dotarray[107][225], dotarray[108][225], dotarray[109][225], dotarray[110][225], dotarray[111][225], dotarray[112][225], dotarray[113][225], dotarray[114][225], dotarray[115][225], dotarray[116][225], dotarray[117][225], dotarray[118][225], dotarray[119][225], dotarray[120][225], dotarray[121][225], dotarray[122][225], dotarray[123][225], dotarray[124][225], dotarray[125][225], dotarray[126][225], dotarray[127][225]};
assign dot_col_226 = {dotarray[0][226], dotarray[1][226], dotarray[2][226], dotarray[3][226], dotarray[4][226], dotarray[5][226], dotarray[6][226], dotarray[7][226], dotarray[8][226], dotarray[9][226], dotarray[10][226], dotarray[11][226], dotarray[12][226], dotarray[13][226], dotarray[14][226], dotarray[15][226], dotarray[16][226], dotarray[17][226], dotarray[18][226], dotarray[19][226], dotarray[20][226], dotarray[21][226], dotarray[22][226], dotarray[23][226], dotarray[24][226], dotarray[25][226], dotarray[26][226], dotarray[27][226], dotarray[28][226], dotarray[29][226], dotarray[30][226], dotarray[31][226], dotarray[32][226], dotarray[33][226], dotarray[34][226], dotarray[35][226], dotarray[36][226], dotarray[37][226], dotarray[38][226], dotarray[39][226], dotarray[40][226], dotarray[41][226], dotarray[42][226], dotarray[43][226], dotarray[44][226], dotarray[45][226], dotarray[46][226], dotarray[47][226], dotarray[48][226], dotarray[49][226], dotarray[50][226], dotarray[51][226], dotarray[52][226], dotarray[53][226], dotarray[54][226], dotarray[55][226], dotarray[56][226], dotarray[57][226], dotarray[58][226], dotarray[59][226], dotarray[60][226], dotarray[61][226], dotarray[62][226], dotarray[63][226], dotarray[64][226], dotarray[65][226], dotarray[66][226], dotarray[67][226], dotarray[68][226], dotarray[69][226], dotarray[70][226], dotarray[71][226], dotarray[72][226], dotarray[73][226], dotarray[74][226], dotarray[75][226], dotarray[76][226], dotarray[77][226], dotarray[78][226], dotarray[79][226], dotarray[80][226], dotarray[81][226], dotarray[82][226], dotarray[83][226], dotarray[84][226], dotarray[85][226], dotarray[86][226], dotarray[87][226], dotarray[88][226], dotarray[89][226], dotarray[90][226], dotarray[91][226], dotarray[92][226], dotarray[93][226], dotarray[94][226], dotarray[95][226], dotarray[96][226], dotarray[97][226], dotarray[98][226], dotarray[99][226], dotarray[100][226], dotarray[101][226], dotarray[102][226], dotarray[103][226], dotarray[104][226], dotarray[105][226], dotarray[106][226], dotarray[107][226], dotarray[108][226], dotarray[109][226], dotarray[110][226], dotarray[111][226], dotarray[112][226], dotarray[113][226], dotarray[114][226], dotarray[115][226], dotarray[116][226], dotarray[117][226], dotarray[118][226], dotarray[119][226], dotarray[120][226], dotarray[121][226], dotarray[122][226], dotarray[123][226], dotarray[124][226], dotarray[125][226], dotarray[126][226], dotarray[127][226]};
assign dot_col_227 = {dotarray[0][227], dotarray[1][227], dotarray[2][227], dotarray[3][227], dotarray[4][227], dotarray[5][227], dotarray[6][227], dotarray[7][227], dotarray[8][227], dotarray[9][227], dotarray[10][227], dotarray[11][227], dotarray[12][227], dotarray[13][227], dotarray[14][227], dotarray[15][227], dotarray[16][227], dotarray[17][227], dotarray[18][227], dotarray[19][227], dotarray[20][227], dotarray[21][227], dotarray[22][227], dotarray[23][227], dotarray[24][227], dotarray[25][227], dotarray[26][227], dotarray[27][227], dotarray[28][227], dotarray[29][227], dotarray[30][227], dotarray[31][227], dotarray[32][227], dotarray[33][227], dotarray[34][227], dotarray[35][227], dotarray[36][227], dotarray[37][227], dotarray[38][227], dotarray[39][227], dotarray[40][227], dotarray[41][227], dotarray[42][227], dotarray[43][227], dotarray[44][227], dotarray[45][227], dotarray[46][227], dotarray[47][227], dotarray[48][227], dotarray[49][227], dotarray[50][227], dotarray[51][227], dotarray[52][227], dotarray[53][227], dotarray[54][227], dotarray[55][227], dotarray[56][227], dotarray[57][227], dotarray[58][227], dotarray[59][227], dotarray[60][227], dotarray[61][227], dotarray[62][227], dotarray[63][227], dotarray[64][227], dotarray[65][227], dotarray[66][227], dotarray[67][227], dotarray[68][227], dotarray[69][227], dotarray[70][227], dotarray[71][227], dotarray[72][227], dotarray[73][227], dotarray[74][227], dotarray[75][227], dotarray[76][227], dotarray[77][227], dotarray[78][227], dotarray[79][227], dotarray[80][227], dotarray[81][227], dotarray[82][227], dotarray[83][227], dotarray[84][227], dotarray[85][227], dotarray[86][227], dotarray[87][227], dotarray[88][227], dotarray[89][227], dotarray[90][227], dotarray[91][227], dotarray[92][227], dotarray[93][227], dotarray[94][227], dotarray[95][227], dotarray[96][227], dotarray[97][227], dotarray[98][227], dotarray[99][227], dotarray[100][227], dotarray[101][227], dotarray[102][227], dotarray[103][227], dotarray[104][227], dotarray[105][227], dotarray[106][227], dotarray[107][227], dotarray[108][227], dotarray[109][227], dotarray[110][227], dotarray[111][227], dotarray[112][227], dotarray[113][227], dotarray[114][227], dotarray[115][227], dotarray[116][227], dotarray[117][227], dotarray[118][227], dotarray[119][227], dotarray[120][227], dotarray[121][227], dotarray[122][227], dotarray[123][227], dotarray[124][227], dotarray[125][227], dotarray[126][227], dotarray[127][227]};
assign dot_col_228 = {dotarray[0][228], dotarray[1][228], dotarray[2][228], dotarray[3][228], dotarray[4][228], dotarray[5][228], dotarray[6][228], dotarray[7][228], dotarray[8][228], dotarray[9][228], dotarray[10][228], dotarray[11][228], dotarray[12][228], dotarray[13][228], dotarray[14][228], dotarray[15][228], dotarray[16][228], dotarray[17][228], dotarray[18][228], dotarray[19][228], dotarray[20][228], dotarray[21][228], dotarray[22][228], dotarray[23][228], dotarray[24][228], dotarray[25][228], dotarray[26][228], dotarray[27][228], dotarray[28][228], dotarray[29][228], dotarray[30][228], dotarray[31][228], dotarray[32][228], dotarray[33][228], dotarray[34][228], dotarray[35][228], dotarray[36][228], dotarray[37][228], dotarray[38][228], dotarray[39][228], dotarray[40][228], dotarray[41][228], dotarray[42][228], dotarray[43][228], dotarray[44][228], dotarray[45][228], dotarray[46][228], dotarray[47][228], dotarray[48][228], dotarray[49][228], dotarray[50][228], dotarray[51][228], dotarray[52][228], dotarray[53][228], dotarray[54][228], dotarray[55][228], dotarray[56][228], dotarray[57][228], dotarray[58][228], dotarray[59][228], dotarray[60][228], dotarray[61][228], dotarray[62][228], dotarray[63][228], dotarray[64][228], dotarray[65][228], dotarray[66][228], dotarray[67][228], dotarray[68][228], dotarray[69][228], dotarray[70][228], dotarray[71][228], dotarray[72][228], dotarray[73][228], dotarray[74][228], dotarray[75][228], dotarray[76][228], dotarray[77][228], dotarray[78][228], dotarray[79][228], dotarray[80][228], dotarray[81][228], dotarray[82][228], dotarray[83][228], dotarray[84][228], dotarray[85][228], dotarray[86][228], dotarray[87][228], dotarray[88][228], dotarray[89][228], dotarray[90][228], dotarray[91][228], dotarray[92][228], dotarray[93][228], dotarray[94][228], dotarray[95][228], dotarray[96][228], dotarray[97][228], dotarray[98][228], dotarray[99][228], dotarray[100][228], dotarray[101][228], dotarray[102][228], dotarray[103][228], dotarray[104][228], dotarray[105][228], dotarray[106][228], dotarray[107][228], dotarray[108][228], dotarray[109][228], dotarray[110][228], dotarray[111][228], dotarray[112][228], dotarray[113][228], dotarray[114][228], dotarray[115][228], dotarray[116][228], dotarray[117][228], dotarray[118][228], dotarray[119][228], dotarray[120][228], dotarray[121][228], dotarray[122][228], dotarray[123][228], dotarray[124][228], dotarray[125][228], dotarray[126][228], dotarray[127][228]};
assign dot_col_229 = {dotarray[0][229], dotarray[1][229], dotarray[2][229], dotarray[3][229], dotarray[4][229], dotarray[5][229], dotarray[6][229], dotarray[7][229], dotarray[8][229], dotarray[9][229], dotarray[10][229], dotarray[11][229], dotarray[12][229], dotarray[13][229], dotarray[14][229], dotarray[15][229], dotarray[16][229], dotarray[17][229], dotarray[18][229], dotarray[19][229], dotarray[20][229], dotarray[21][229], dotarray[22][229], dotarray[23][229], dotarray[24][229], dotarray[25][229], dotarray[26][229], dotarray[27][229], dotarray[28][229], dotarray[29][229], dotarray[30][229], dotarray[31][229], dotarray[32][229], dotarray[33][229], dotarray[34][229], dotarray[35][229], dotarray[36][229], dotarray[37][229], dotarray[38][229], dotarray[39][229], dotarray[40][229], dotarray[41][229], dotarray[42][229], dotarray[43][229], dotarray[44][229], dotarray[45][229], dotarray[46][229], dotarray[47][229], dotarray[48][229], dotarray[49][229], dotarray[50][229], dotarray[51][229], dotarray[52][229], dotarray[53][229], dotarray[54][229], dotarray[55][229], dotarray[56][229], dotarray[57][229], dotarray[58][229], dotarray[59][229], dotarray[60][229], dotarray[61][229], dotarray[62][229], dotarray[63][229], dotarray[64][229], dotarray[65][229], dotarray[66][229], dotarray[67][229], dotarray[68][229], dotarray[69][229], dotarray[70][229], dotarray[71][229], dotarray[72][229], dotarray[73][229], dotarray[74][229], dotarray[75][229], dotarray[76][229], dotarray[77][229], dotarray[78][229], dotarray[79][229], dotarray[80][229], dotarray[81][229], dotarray[82][229], dotarray[83][229], dotarray[84][229], dotarray[85][229], dotarray[86][229], dotarray[87][229], dotarray[88][229], dotarray[89][229], dotarray[90][229], dotarray[91][229], dotarray[92][229], dotarray[93][229], dotarray[94][229], dotarray[95][229], dotarray[96][229], dotarray[97][229], dotarray[98][229], dotarray[99][229], dotarray[100][229], dotarray[101][229], dotarray[102][229], dotarray[103][229], dotarray[104][229], dotarray[105][229], dotarray[106][229], dotarray[107][229], dotarray[108][229], dotarray[109][229], dotarray[110][229], dotarray[111][229], dotarray[112][229], dotarray[113][229], dotarray[114][229], dotarray[115][229], dotarray[116][229], dotarray[117][229], dotarray[118][229], dotarray[119][229], dotarray[120][229], dotarray[121][229], dotarray[122][229], dotarray[123][229], dotarray[124][229], dotarray[125][229], dotarray[126][229], dotarray[127][229]};
assign dot_col_230 = {dotarray[0][230], dotarray[1][230], dotarray[2][230], dotarray[3][230], dotarray[4][230], dotarray[5][230], dotarray[6][230], dotarray[7][230], dotarray[8][230], dotarray[9][230], dotarray[10][230], dotarray[11][230], dotarray[12][230], dotarray[13][230], dotarray[14][230], dotarray[15][230], dotarray[16][230], dotarray[17][230], dotarray[18][230], dotarray[19][230], dotarray[20][230], dotarray[21][230], dotarray[22][230], dotarray[23][230], dotarray[24][230], dotarray[25][230], dotarray[26][230], dotarray[27][230], dotarray[28][230], dotarray[29][230], dotarray[30][230], dotarray[31][230], dotarray[32][230], dotarray[33][230], dotarray[34][230], dotarray[35][230], dotarray[36][230], dotarray[37][230], dotarray[38][230], dotarray[39][230], dotarray[40][230], dotarray[41][230], dotarray[42][230], dotarray[43][230], dotarray[44][230], dotarray[45][230], dotarray[46][230], dotarray[47][230], dotarray[48][230], dotarray[49][230], dotarray[50][230], dotarray[51][230], dotarray[52][230], dotarray[53][230], dotarray[54][230], dotarray[55][230], dotarray[56][230], dotarray[57][230], dotarray[58][230], dotarray[59][230], dotarray[60][230], dotarray[61][230], dotarray[62][230], dotarray[63][230], dotarray[64][230], dotarray[65][230], dotarray[66][230], dotarray[67][230], dotarray[68][230], dotarray[69][230], dotarray[70][230], dotarray[71][230], dotarray[72][230], dotarray[73][230], dotarray[74][230], dotarray[75][230], dotarray[76][230], dotarray[77][230], dotarray[78][230], dotarray[79][230], dotarray[80][230], dotarray[81][230], dotarray[82][230], dotarray[83][230], dotarray[84][230], dotarray[85][230], dotarray[86][230], dotarray[87][230], dotarray[88][230], dotarray[89][230], dotarray[90][230], dotarray[91][230], dotarray[92][230], dotarray[93][230], dotarray[94][230], dotarray[95][230], dotarray[96][230], dotarray[97][230], dotarray[98][230], dotarray[99][230], dotarray[100][230], dotarray[101][230], dotarray[102][230], dotarray[103][230], dotarray[104][230], dotarray[105][230], dotarray[106][230], dotarray[107][230], dotarray[108][230], dotarray[109][230], dotarray[110][230], dotarray[111][230], dotarray[112][230], dotarray[113][230], dotarray[114][230], dotarray[115][230], dotarray[116][230], dotarray[117][230], dotarray[118][230], dotarray[119][230], dotarray[120][230], dotarray[121][230], dotarray[122][230], dotarray[123][230], dotarray[124][230], dotarray[125][230], dotarray[126][230], dotarray[127][230]};
assign dot_col_231 = {dotarray[0][231], dotarray[1][231], dotarray[2][231], dotarray[3][231], dotarray[4][231], dotarray[5][231], dotarray[6][231], dotarray[7][231], dotarray[8][231], dotarray[9][231], dotarray[10][231], dotarray[11][231], dotarray[12][231], dotarray[13][231], dotarray[14][231], dotarray[15][231], dotarray[16][231], dotarray[17][231], dotarray[18][231], dotarray[19][231], dotarray[20][231], dotarray[21][231], dotarray[22][231], dotarray[23][231], dotarray[24][231], dotarray[25][231], dotarray[26][231], dotarray[27][231], dotarray[28][231], dotarray[29][231], dotarray[30][231], dotarray[31][231], dotarray[32][231], dotarray[33][231], dotarray[34][231], dotarray[35][231], dotarray[36][231], dotarray[37][231], dotarray[38][231], dotarray[39][231], dotarray[40][231], dotarray[41][231], dotarray[42][231], dotarray[43][231], dotarray[44][231], dotarray[45][231], dotarray[46][231], dotarray[47][231], dotarray[48][231], dotarray[49][231], dotarray[50][231], dotarray[51][231], dotarray[52][231], dotarray[53][231], dotarray[54][231], dotarray[55][231], dotarray[56][231], dotarray[57][231], dotarray[58][231], dotarray[59][231], dotarray[60][231], dotarray[61][231], dotarray[62][231], dotarray[63][231], dotarray[64][231], dotarray[65][231], dotarray[66][231], dotarray[67][231], dotarray[68][231], dotarray[69][231], dotarray[70][231], dotarray[71][231], dotarray[72][231], dotarray[73][231], dotarray[74][231], dotarray[75][231], dotarray[76][231], dotarray[77][231], dotarray[78][231], dotarray[79][231], dotarray[80][231], dotarray[81][231], dotarray[82][231], dotarray[83][231], dotarray[84][231], dotarray[85][231], dotarray[86][231], dotarray[87][231], dotarray[88][231], dotarray[89][231], dotarray[90][231], dotarray[91][231], dotarray[92][231], dotarray[93][231], dotarray[94][231], dotarray[95][231], dotarray[96][231], dotarray[97][231], dotarray[98][231], dotarray[99][231], dotarray[100][231], dotarray[101][231], dotarray[102][231], dotarray[103][231], dotarray[104][231], dotarray[105][231], dotarray[106][231], dotarray[107][231], dotarray[108][231], dotarray[109][231], dotarray[110][231], dotarray[111][231], dotarray[112][231], dotarray[113][231], dotarray[114][231], dotarray[115][231], dotarray[116][231], dotarray[117][231], dotarray[118][231], dotarray[119][231], dotarray[120][231], dotarray[121][231], dotarray[122][231], dotarray[123][231], dotarray[124][231], dotarray[125][231], dotarray[126][231], dotarray[127][231]};
assign dot_col_232 = {dotarray[0][232], dotarray[1][232], dotarray[2][232], dotarray[3][232], dotarray[4][232], dotarray[5][232], dotarray[6][232], dotarray[7][232], dotarray[8][232], dotarray[9][232], dotarray[10][232], dotarray[11][232], dotarray[12][232], dotarray[13][232], dotarray[14][232], dotarray[15][232], dotarray[16][232], dotarray[17][232], dotarray[18][232], dotarray[19][232], dotarray[20][232], dotarray[21][232], dotarray[22][232], dotarray[23][232], dotarray[24][232], dotarray[25][232], dotarray[26][232], dotarray[27][232], dotarray[28][232], dotarray[29][232], dotarray[30][232], dotarray[31][232], dotarray[32][232], dotarray[33][232], dotarray[34][232], dotarray[35][232], dotarray[36][232], dotarray[37][232], dotarray[38][232], dotarray[39][232], dotarray[40][232], dotarray[41][232], dotarray[42][232], dotarray[43][232], dotarray[44][232], dotarray[45][232], dotarray[46][232], dotarray[47][232], dotarray[48][232], dotarray[49][232], dotarray[50][232], dotarray[51][232], dotarray[52][232], dotarray[53][232], dotarray[54][232], dotarray[55][232], dotarray[56][232], dotarray[57][232], dotarray[58][232], dotarray[59][232], dotarray[60][232], dotarray[61][232], dotarray[62][232], dotarray[63][232], dotarray[64][232], dotarray[65][232], dotarray[66][232], dotarray[67][232], dotarray[68][232], dotarray[69][232], dotarray[70][232], dotarray[71][232], dotarray[72][232], dotarray[73][232], dotarray[74][232], dotarray[75][232], dotarray[76][232], dotarray[77][232], dotarray[78][232], dotarray[79][232], dotarray[80][232], dotarray[81][232], dotarray[82][232], dotarray[83][232], dotarray[84][232], dotarray[85][232], dotarray[86][232], dotarray[87][232], dotarray[88][232], dotarray[89][232], dotarray[90][232], dotarray[91][232], dotarray[92][232], dotarray[93][232], dotarray[94][232], dotarray[95][232], dotarray[96][232], dotarray[97][232], dotarray[98][232], dotarray[99][232], dotarray[100][232], dotarray[101][232], dotarray[102][232], dotarray[103][232], dotarray[104][232], dotarray[105][232], dotarray[106][232], dotarray[107][232], dotarray[108][232], dotarray[109][232], dotarray[110][232], dotarray[111][232], dotarray[112][232], dotarray[113][232], dotarray[114][232], dotarray[115][232], dotarray[116][232], dotarray[117][232], dotarray[118][232], dotarray[119][232], dotarray[120][232], dotarray[121][232], dotarray[122][232], dotarray[123][232], dotarray[124][232], dotarray[125][232], dotarray[126][232], dotarray[127][232]};
assign dot_col_233 = {dotarray[0][233], dotarray[1][233], dotarray[2][233], dotarray[3][233], dotarray[4][233], dotarray[5][233], dotarray[6][233], dotarray[7][233], dotarray[8][233], dotarray[9][233], dotarray[10][233], dotarray[11][233], dotarray[12][233], dotarray[13][233], dotarray[14][233], dotarray[15][233], dotarray[16][233], dotarray[17][233], dotarray[18][233], dotarray[19][233], dotarray[20][233], dotarray[21][233], dotarray[22][233], dotarray[23][233], dotarray[24][233], dotarray[25][233], dotarray[26][233], dotarray[27][233], dotarray[28][233], dotarray[29][233], dotarray[30][233], dotarray[31][233], dotarray[32][233], dotarray[33][233], dotarray[34][233], dotarray[35][233], dotarray[36][233], dotarray[37][233], dotarray[38][233], dotarray[39][233], dotarray[40][233], dotarray[41][233], dotarray[42][233], dotarray[43][233], dotarray[44][233], dotarray[45][233], dotarray[46][233], dotarray[47][233], dotarray[48][233], dotarray[49][233], dotarray[50][233], dotarray[51][233], dotarray[52][233], dotarray[53][233], dotarray[54][233], dotarray[55][233], dotarray[56][233], dotarray[57][233], dotarray[58][233], dotarray[59][233], dotarray[60][233], dotarray[61][233], dotarray[62][233], dotarray[63][233], dotarray[64][233], dotarray[65][233], dotarray[66][233], dotarray[67][233], dotarray[68][233], dotarray[69][233], dotarray[70][233], dotarray[71][233], dotarray[72][233], dotarray[73][233], dotarray[74][233], dotarray[75][233], dotarray[76][233], dotarray[77][233], dotarray[78][233], dotarray[79][233], dotarray[80][233], dotarray[81][233], dotarray[82][233], dotarray[83][233], dotarray[84][233], dotarray[85][233], dotarray[86][233], dotarray[87][233], dotarray[88][233], dotarray[89][233], dotarray[90][233], dotarray[91][233], dotarray[92][233], dotarray[93][233], dotarray[94][233], dotarray[95][233], dotarray[96][233], dotarray[97][233], dotarray[98][233], dotarray[99][233], dotarray[100][233], dotarray[101][233], dotarray[102][233], dotarray[103][233], dotarray[104][233], dotarray[105][233], dotarray[106][233], dotarray[107][233], dotarray[108][233], dotarray[109][233], dotarray[110][233], dotarray[111][233], dotarray[112][233], dotarray[113][233], dotarray[114][233], dotarray[115][233], dotarray[116][233], dotarray[117][233], dotarray[118][233], dotarray[119][233], dotarray[120][233], dotarray[121][233], dotarray[122][233], dotarray[123][233], dotarray[124][233], dotarray[125][233], dotarray[126][233], dotarray[127][233]};
assign dot_col_234 = {dotarray[0][234], dotarray[1][234], dotarray[2][234], dotarray[3][234], dotarray[4][234], dotarray[5][234], dotarray[6][234], dotarray[7][234], dotarray[8][234], dotarray[9][234], dotarray[10][234], dotarray[11][234], dotarray[12][234], dotarray[13][234], dotarray[14][234], dotarray[15][234], dotarray[16][234], dotarray[17][234], dotarray[18][234], dotarray[19][234], dotarray[20][234], dotarray[21][234], dotarray[22][234], dotarray[23][234], dotarray[24][234], dotarray[25][234], dotarray[26][234], dotarray[27][234], dotarray[28][234], dotarray[29][234], dotarray[30][234], dotarray[31][234], dotarray[32][234], dotarray[33][234], dotarray[34][234], dotarray[35][234], dotarray[36][234], dotarray[37][234], dotarray[38][234], dotarray[39][234], dotarray[40][234], dotarray[41][234], dotarray[42][234], dotarray[43][234], dotarray[44][234], dotarray[45][234], dotarray[46][234], dotarray[47][234], dotarray[48][234], dotarray[49][234], dotarray[50][234], dotarray[51][234], dotarray[52][234], dotarray[53][234], dotarray[54][234], dotarray[55][234], dotarray[56][234], dotarray[57][234], dotarray[58][234], dotarray[59][234], dotarray[60][234], dotarray[61][234], dotarray[62][234], dotarray[63][234], dotarray[64][234], dotarray[65][234], dotarray[66][234], dotarray[67][234], dotarray[68][234], dotarray[69][234], dotarray[70][234], dotarray[71][234], dotarray[72][234], dotarray[73][234], dotarray[74][234], dotarray[75][234], dotarray[76][234], dotarray[77][234], dotarray[78][234], dotarray[79][234], dotarray[80][234], dotarray[81][234], dotarray[82][234], dotarray[83][234], dotarray[84][234], dotarray[85][234], dotarray[86][234], dotarray[87][234], dotarray[88][234], dotarray[89][234], dotarray[90][234], dotarray[91][234], dotarray[92][234], dotarray[93][234], dotarray[94][234], dotarray[95][234], dotarray[96][234], dotarray[97][234], dotarray[98][234], dotarray[99][234], dotarray[100][234], dotarray[101][234], dotarray[102][234], dotarray[103][234], dotarray[104][234], dotarray[105][234], dotarray[106][234], dotarray[107][234], dotarray[108][234], dotarray[109][234], dotarray[110][234], dotarray[111][234], dotarray[112][234], dotarray[113][234], dotarray[114][234], dotarray[115][234], dotarray[116][234], dotarray[117][234], dotarray[118][234], dotarray[119][234], dotarray[120][234], dotarray[121][234], dotarray[122][234], dotarray[123][234], dotarray[124][234], dotarray[125][234], dotarray[126][234], dotarray[127][234]};
assign dot_col_235 = {dotarray[0][235], dotarray[1][235], dotarray[2][235], dotarray[3][235], dotarray[4][235], dotarray[5][235], dotarray[6][235], dotarray[7][235], dotarray[8][235], dotarray[9][235], dotarray[10][235], dotarray[11][235], dotarray[12][235], dotarray[13][235], dotarray[14][235], dotarray[15][235], dotarray[16][235], dotarray[17][235], dotarray[18][235], dotarray[19][235], dotarray[20][235], dotarray[21][235], dotarray[22][235], dotarray[23][235], dotarray[24][235], dotarray[25][235], dotarray[26][235], dotarray[27][235], dotarray[28][235], dotarray[29][235], dotarray[30][235], dotarray[31][235], dotarray[32][235], dotarray[33][235], dotarray[34][235], dotarray[35][235], dotarray[36][235], dotarray[37][235], dotarray[38][235], dotarray[39][235], dotarray[40][235], dotarray[41][235], dotarray[42][235], dotarray[43][235], dotarray[44][235], dotarray[45][235], dotarray[46][235], dotarray[47][235], dotarray[48][235], dotarray[49][235], dotarray[50][235], dotarray[51][235], dotarray[52][235], dotarray[53][235], dotarray[54][235], dotarray[55][235], dotarray[56][235], dotarray[57][235], dotarray[58][235], dotarray[59][235], dotarray[60][235], dotarray[61][235], dotarray[62][235], dotarray[63][235], dotarray[64][235], dotarray[65][235], dotarray[66][235], dotarray[67][235], dotarray[68][235], dotarray[69][235], dotarray[70][235], dotarray[71][235], dotarray[72][235], dotarray[73][235], dotarray[74][235], dotarray[75][235], dotarray[76][235], dotarray[77][235], dotarray[78][235], dotarray[79][235], dotarray[80][235], dotarray[81][235], dotarray[82][235], dotarray[83][235], dotarray[84][235], dotarray[85][235], dotarray[86][235], dotarray[87][235], dotarray[88][235], dotarray[89][235], dotarray[90][235], dotarray[91][235], dotarray[92][235], dotarray[93][235], dotarray[94][235], dotarray[95][235], dotarray[96][235], dotarray[97][235], dotarray[98][235], dotarray[99][235], dotarray[100][235], dotarray[101][235], dotarray[102][235], dotarray[103][235], dotarray[104][235], dotarray[105][235], dotarray[106][235], dotarray[107][235], dotarray[108][235], dotarray[109][235], dotarray[110][235], dotarray[111][235], dotarray[112][235], dotarray[113][235], dotarray[114][235], dotarray[115][235], dotarray[116][235], dotarray[117][235], dotarray[118][235], dotarray[119][235], dotarray[120][235], dotarray[121][235], dotarray[122][235], dotarray[123][235], dotarray[124][235], dotarray[125][235], dotarray[126][235], dotarray[127][235]};
assign dot_col_236 = {dotarray[0][236], dotarray[1][236], dotarray[2][236], dotarray[3][236], dotarray[4][236], dotarray[5][236], dotarray[6][236], dotarray[7][236], dotarray[8][236], dotarray[9][236], dotarray[10][236], dotarray[11][236], dotarray[12][236], dotarray[13][236], dotarray[14][236], dotarray[15][236], dotarray[16][236], dotarray[17][236], dotarray[18][236], dotarray[19][236], dotarray[20][236], dotarray[21][236], dotarray[22][236], dotarray[23][236], dotarray[24][236], dotarray[25][236], dotarray[26][236], dotarray[27][236], dotarray[28][236], dotarray[29][236], dotarray[30][236], dotarray[31][236], dotarray[32][236], dotarray[33][236], dotarray[34][236], dotarray[35][236], dotarray[36][236], dotarray[37][236], dotarray[38][236], dotarray[39][236], dotarray[40][236], dotarray[41][236], dotarray[42][236], dotarray[43][236], dotarray[44][236], dotarray[45][236], dotarray[46][236], dotarray[47][236], dotarray[48][236], dotarray[49][236], dotarray[50][236], dotarray[51][236], dotarray[52][236], dotarray[53][236], dotarray[54][236], dotarray[55][236], dotarray[56][236], dotarray[57][236], dotarray[58][236], dotarray[59][236], dotarray[60][236], dotarray[61][236], dotarray[62][236], dotarray[63][236], dotarray[64][236], dotarray[65][236], dotarray[66][236], dotarray[67][236], dotarray[68][236], dotarray[69][236], dotarray[70][236], dotarray[71][236], dotarray[72][236], dotarray[73][236], dotarray[74][236], dotarray[75][236], dotarray[76][236], dotarray[77][236], dotarray[78][236], dotarray[79][236], dotarray[80][236], dotarray[81][236], dotarray[82][236], dotarray[83][236], dotarray[84][236], dotarray[85][236], dotarray[86][236], dotarray[87][236], dotarray[88][236], dotarray[89][236], dotarray[90][236], dotarray[91][236], dotarray[92][236], dotarray[93][236], dotarray[94][236], dotarray[95][236], dotarray[96][236], dotarray[97][236], dotarray[98][236], dotarray[99][236], dotarray[100][236], dotarray[101][236], dotarray[102][236], dotarray[103][236], dotarray[104][236], dotarray[105][236], dotarray[106][236], dotarray[107][236], dotarray[108][236], dotarray[109][236], dotarray[110][236], dotarray[111][236], dotarray[112][236], dotarray[113][236], dotarray[114][236], dotarray[115][236], dotarray[116][236], dotarray[117][236], dotarray[118][236], dotarray[119][236], dotarray[120][236], dotarray[121][236], dotarray[122][236], dotarray[123][236], dotarray[124][236], dotarray[125][236], dotarray[126][236], dotarray[127][236]};
assign dot_col_237 = {dotarray[0][237], dotarray[1][237], dotarray[2][237], dotarray[3][237], dotarray[4][237], dotarray[5][237], dotarray[6][237], dotarray[7][237], dotarray[8][237], dotarray[9][237], dotarray[10][237], dotarray[11][237], dotarray[12][237], dotarray[13][237], dotarray[14][237], dotarray[15][237], dotarray[16][237], dotarray[17][237], dotarray[18][237], dotarray[19][237], dotarray[20][237], dotarray[21][237], dotarray[22][237], dotarray[23][237], dotarray[24][237], dotarray[25][237], dotarray[26][237], dotarray[27][237], dotarray[28][237], dotarray[29][237], dotarray[30][237], dotarray[31][237], dotarray[32][237], dotarray[33][237], dotarray[34][237], dotarray[35][237], dotarray[36][237], dotarray[37][237], dotarray[38][237], dotarray[39][237], dotarray[40][237], dotarray[41][237], dotarray[42][237], dotarray[43][237], dotarray[44][237], dotarray[45][237], dotarray[46][237], dotarray[47][237], dotarray[48][237], dotarray[49][237], dotarray[50][237], dotarray[51][237], dotarray[52][237], dotarray[53][237], dotarray[54][237], dotarray[55][237], dotarray[56][237], dotarray[57][237], dotarray[58][237], dotarray[59][237], dotarray[60][237], dotarray[61][237], dotarray[62][237], dotarray[63][237], dotarray[64][237], dotarray[65][237], dotarray[66][237], dotarray[67][237], dotarray[68][237], dotarray[69][237], dotarray[70][237], dotarray[71][237], dotarray[72][237], dotarray[73][237], dotarray[74][237], dotarray[75][237], dotarray[76][237], dotarray[77][237], dotarray[78][237], dotarray[79][237], dotarray[80][237], dotarray[81][237], dotarray[82][237], dotarray[83][237], dotarray[84][237], dotarray[85][237], dotarray[86][237], dotarray[87][237], dotarray[88][237], dotarray[89][237], dotarray[90][237], dotarray[91][237], dotarray[92][237], dotarray[93][237], dotarray[94][237], dotarray[95][237], dotarray[96][237], dotarray[97][237], dotarray[98][237], dotarray[99][237], dotarray[100][237], dotarray[101][237], dotarray[102][237], dotarray[103][237], dotarray[104][237], dotarray[105][237], dotarray[106][237], dotarray[107][237], dotarray[108][237], dotarray[109][237], dotarray[110][237], dotarray[111][237], dotarray[112][237], dotarray[113][237], dotarray[114][237], dotarray[115][237], dotarray[116][237], dotarray[117][237], dotarray[118][237], dotarray[119][237], dotarray[120][237], dotarray[121][237], dotarray[122][237], dotarray[123][237], dotarray[124][237], dotarray[125][237], dotarray[126][237], dotarray[127][237]};
assign dot_col_238 = {dotarray[0][238], dotarray[1][238], dotarray[2][238], dotarray[3][238], dotarray[4][238], dotarray[5][238], dotarray[6][238], dotarray[7][238], dotarray[8][238], dotarray[9][238], dotarray[10][238], dotarray[11][238], dotarray[12][238], dotarray[13][238], dotarray[14][238], dotarray[15][238], dotarray[16][238], dotarray[17][238], dotarray[18][238], dotarray[19][238], dotarray[20][238], dotarray[21][238], dotarray[22][238], dotarray[23][238], dotarray[24][238], dotarray[25][238], dotarray[26][238], dotarray[27][238], dotarray[28][238], dotarray[29][238], dotarray[30][238], dotarray[31][238], dotarray[32][238], dotarray[33][238], dotarray[34][238], dotarray[35][238], dotarray[36][238], dotarray[37][238], dotarray[38][238], dotarray[39][238], dotarray[40][238], dotarray[41][238], dotarray[42][238], dotarray[43][238], dotarray[44][238], dotarray[45][238], dotarray[46][238], dotarray[47][238], dotarray[48][238], dotarray[49][238], dotarray[50][238], dotarray[51][238], dotarray[52][238], dotarray[53][238], dotarray[54][238], dotarray[55][238], dotarray[56][238], dotarray[57][238], dotarray[58][238], dotarray[59][238], dotarray[60][238], dotarray[61][238], dotarray[62][238], dotarray[63][238], dotarray[64][238], dotarray[65][238], dotarray[66][238], dotarray[67][238], dotarray[68][238], dotarray[69][238], dotarray[70][238], dotarray[71][238], dotarray[72][238], dotarray[73][238], dotarray[74][238], dotarray[75][238], dotarray[76][238], dotarray[77][238], dotarray[78][238], dotarray[79][238], dotarray[80][238], dotarray[81][238], dotarray[82][238], dotarray[83][238], dotarray[84][238], dotarray[85][238], dotarray[86][238], dotarray[87][238], dotarray[88][238], dotarray[89][238], dotarray[90][238], dotarray[91][238], dotarray[92][238], dotarray[93][238], dotarray[94][238], dotarray[95][238], dotarray[96][238], dotarray[97][238], dotarray[98][238], dotarray[99][238], dotarray[100][238], dotarray[101][238], dotarray[102][238], dotarray[103][238], dotarray[104][238], dotarray[105][238], dotarray[106][238], dotarray[107][238], dotarray[108][238], dotarray[109][238], dotarray[110][238], dotarray[111][238], dotarray[112][238], dotarray[113][238], dotarray[114][238], dotarray[115][238], dotarray[116][238], dotarray[117][238], dotarray[118][238], dotarray[119][238], dotarray[120][238], dotarray[121][238], dotarray[122][238], dotarray[123][238], dotarray[124][238], dotarray[125][238], dotarray[126][238], dotarray[127][238]};
assign dot_col_239 = {dotarray[0][239], dotarray[1][239], dotarray[2][239], dotarray[3][239], dotarray[4][239], dotarray[5][239], dotarray[6][239], dotarray[7][239], dotarray[8][239], dotarray[9][239], dotarray[10][239], dotarray[11][239], dotarray[12][239], dotarray[13][239], dotarray[14][239], dotarray[15][239], dotarray[16][239], dotarray[17][239], dotarray[18][239], dotarray[19][239], dotarray[20][239], dotarray[21][239], dotarray[22][239], dotarray[23][239], dotarray[24][239], dotarray[25][239], dotarray[26][239], dotarray[27][239], dotarray[28][239], dotarray[29][239], dotarray[30][239], dotarray[31][239], dotarray[32][239], dotarray[33][239], dotarray[34][239], dotarray[35][239], dotarray[36][239], dotarray[37][239], dotarray[38][239], dotarray[39][239], dotarray[40][239], dotarray[41][239], dotarray[42][239], dotarray[43][239], dotarray[44][239], dotarray[45][239], dotarray[46][239], dotarray[47][239], dotarray[48][239], dotarray[49][239], dotarray[50][239], dotarray[51][239], dotarray[52][239], dotarray[53][239], dotarray[54][239], dotarray[55][239], dotarray[56][239], dotarray[57][239], dotarray[58][239], dotarray[59][239], dotarray[60][239], dotarray[61][239], dotarray[62][239], dotarray[63][239], dotarray[64][239], dotarray[65][239], dotarray[66][239], dotarray[67][239], dotarray[68][239], dotarray[69][239], dotarray[70][239], dotarray[71][239], dotarray[72][239], dotarray[73][239], dotarray[74][239], dotarray[75][239], dotarray[76][239], dotarray[77][239], dotarray[78][239], dotarray[79][239], dotarray[80][239], dotarray[81][239], dotarray[82][239], dotarray[83][239], dotarray[84][239], dotarray[85][239], dotarray[86][239], dotarray[87][239], dotarray[88][239], dotarray[89][239], dotarray[90][239], dotarray[91][239], dotarray[92][239], dotarray[93][239], dotarray[94][239], dotarray[95][239], dotarray[96][239], dotarray[97][239], dotarray[98][239], dotarray[99][239], dotarray[100][239], dotarray[101][239], dotarray[102][239], dotarray[103][239], dotarray[104][239], dotarray[105][239], dotarray[106][239], dotarray[107][239], dotarray[108][239], dotarray[109][239], dotarray[110][239], dotarray[111][239], dotarray[112][239], dotarray[113][239], dotarray[114][239], dotarray[115][239], dotarray[116][239], dotarray[117][239], dotarray[118][239], dotarray[119][239], dotarray[120][239], dotarray[121][239], dotarray[122][239], dotarray[123][239], dotarray[124][239], dotarray[125][239], dotarray[126][239], dotarray[127][239]};
assign dot_col_240 = {dotarray[0][240], dotarray[1][240], dotarray[2][240], dotarray[3][240], dotarray[4][240], dotarray[5][240], dotarray[6][240], dotarray[7][240], dotarray[8][240], dotarray[9][240], dotarray[10][240], dotarray[11][240], dotarray[12][240], dotarray[13][240], dotarray[14][240], dotarray[15][240], dotarray[16][240], dotarray[17][240], dotarray[18][240], dotarray[19][240], dotarray[20][240], dotarray[21][240], dotarray[22][240], dotarray[23][240], dotarray[24][240], dotarray[25][240], dotarray[26][240], dotarray[27][240], dotarray[28][240], dotarray[29][240], dotarray[30][240], dotarray[31][240], dotarray[32][240], dotarray[33][240], dotarray[34][240], dotarray[35][240], dotarray[36][240], dotarray[37][240], dotarray[38][240], dotarray[39][240], dotarray[40][240], dotarray[41][240], dotarray[42][240], dotarray[43][240], dotarray[44][240], dotarray[45][240], dotarray[46][240], dotarray[47][240], dotarray[48][240], dotarray[49][240], dotarray[50][240], dotarray[51][240], dotarray[52][240], dotarray[53][240], dotarray[54][240], dotarray[55][240], dotarray[56][240], dotarray[57][240], dotarray[58][240], dotarray[59][240], dotarray[60][240], dotarray[61][240], dotarray[62][240], dotarray[63][240], dotarray[64][240], dotarray[65][240], dotarray[66][240], dotarray[67][240], dotarray[68][240], dotarray[69][240], dotarray[70][240], dotarray[71][240], dotarray[72][240], dotarray[73][240], dotarray[74][240], dotarray[75][240], dotarray[76][240], dotarray[77][240], dotarray[78][240], dotarray[79][240], dotarray[80][240], dotarray[81][240], dotarray[82][240], dotarray[83][240], dotarray[84][240], dotarray[85][240], dotarray[86][240], dotarray[87][240], dotarray[88][240], dotarray[89][240], dotarray[90][240], dotarray[91][240], dotarray[92][240], dotarray[93][240], dotarray[94][240], dotarray[95][240], dotarray[96][240], dotarray[97][240], dotarray[98][240], dotarray[99][240], dotarray[100][240], dotarray[101][240], dotarray[102][240], dotarray[103][240], dotarray[104][240], dotarray[105][240], dotarray[106][240], dotarray[107][240], dotarray[108][240], dotarray[109][240], dotarray[110][240], dotarray[111][240], dotarray[112][240], dotarray[113][240], dotarray[114][240], dotarray[115][240], dotarray[116][240], dotarray[117][240], dotarray[118][240], dotarray[119][240], dotarray[120][240], dotarray[121][240], dotarray[122][240], dotarray[123][240], dotarray[124][240], dotarray[125][240], dotarray[126][240], dotarray[127][240]};
assign dot_col_241 = {dotarray[0][241], dotarray[1][241], dotarray[2][241], dotarray[3][241], dotarray[4][241], dotarray[5][241], dotarray[6][241], dotarray[7][241], dotarray[8][241], dotarray[9][241], dotarray[10][241], dotarray[11][241], dotarray[12][241], dotarray[13][241], dotarray[14][241], dotarray[15][241], dotarray[16][241], dotarray[17][241], dotarray[18][241], dotarray[19][241], dotarray[20][241], dotarray[21][241], dotarray[22][241], dotarray[23][241], dotarray[24][241], dotarray[25][241], dotarray[26][241], dotarray[27][241], dotarray[28][241], dotarray[29][241], dotarray[30][241], dotarray[31][241], dotarray[32][241], dotarray[33][241], dotarray[34][241], dotarray[35][241], dotarray[36][241], dotarray[37][241], dotarray[38][241], dotarray[39][241], dotarray[40][241], dotarray[41][241], dotarray[42][241], dotarray[43][241], dotarray[44][241], dotarray[45][241], dotarray[46][241], dotarray[47][241], dotarray[48][241], dotarray[49][241], dotarray[50][241], dotarray[51][241], dotarray[52][241], dotarray[53][241], dotarray[54][241], dotarray[55][241], dotarray[56][241], dotarray[57][241], dotarray[58][241], dotarray[59][241], dotarray[60][241], dotarray[61][241], dotarray[62][241], dotarray[63][241], dotarray[64][241], dotarray[65][241], dotarray[66][241], dotarray[67][241], dotarray[68][241], dotarray[69][241], dotarray[70][241], dotarray[71][241], dotarray[72][241], dotarray[73][241], dotarray[74][241], dotarray[75][241], dotarray[76][241], dotarray[77][241], dotarray[78][241], dotarray[79][241], dotarray[80][241], dotarray[81][241], dotarray[82][241], dotarray[83][241], dotarray[84][241], dotarray[85][241], dotarray[86][241], dotarray[87][241], dotarray[88][241], dotarray[89][241], dotarray[90][241], dotarray[91][241], dotarray[92][241], dotarray[93][241], dotarray[94][241], dotarray[95][241], dotarray[96][241], dotarray[97][241], dotarray[98][241], dotarray[99][241], dotarray[100][241], dotarray[101][241], dotarray[102][241], dotarray[103][241], dotarray[104][241], dotarray[105][241], dotarray[106][241], dotarray[107][241], dotarray[108][241], dotarray[109][241], dotarray[110][241], dotarray[111][241], dotarray[112][241], dotarray[113][241], dotarray[114][241], dotarray[115][241], dotarray[116][241], dotarray[117][241], dotarray[118][241], dotarray[119][241], dotarray[120][241], dotarray[121][241], dotarray[122][241], dotarray[123][241], dotarray[124][241], dotarray[125][241], dotarray[126][241], dotarray[127][241]};
assign dot_col_242 = {dotarray[0][242], dotarray[1][242], dotarray[2][242], dotarray[3][242], dotarray[4][242], dotarray[5][242], dotarray[6][242], dotarray[7][242], dotarray[8][242], dotarray[9][242], dotarray[10][242], dotarray[11][242], dotarray[12][242], dotarray[13][242], dotarray[14][242], dotarray[15][242], dotarray[16][242], dotarray[17][242], dotarray[18][242], dotarray[19][242], dotarray[20][242], dotarray[21][242], dotarray[22][242], dotarray[23][242], dotarray[24][242], dotarray[25][242], dotarray[26][242], dotarray[27][242], dotarray[28][242], dotarray[29][242], dotarray[30][242], dotarray[31][242], dotarray[32][242], dotarray[33][242], dotarray[34][242], dotarray[35][242], dotarray[36][242], dotarray[37][242], dotarray[38][242], dotarray[39][242], dotarray[40][242], dotarray[41][242], dotarray[42][242], dotarray[43][242], dotarray[44][242], dotarray[45][242], dotarray[46][242], dotarray[47][242], dotarray[48][242], dotarray[49][242], dotarray[50][242], dotarray[51][242], dotarray[52][242], dotarray[53][242], dotarray[54][242], dotarray[55][242], dotarray[56][242], dotarray[57][242], dotarray[58][242], dotarray[59][242], dotarray[60][242], dotarray[61][242], dotarray[62][242], dotarray[63][242], dotarray[64][242], dotarray[65][242], dotarray[66][242], dotarray[67][242], dotarray[68][242], dotarray[69][242], dotarray[70][242], dotarray[71][242], dotarray[72][242], dotarray[73][242], dotarray[74][242], dotarray[75][242], dotarray[76][242], dotarray[77][242], dotarray[78][242], dotarray[79][242], dotarray[80][242], dotarray[81][242], dotarray[82][242], dotarray[83][242], dotarray[84][242], dotarray[85][242], dotarray[86][242], dotarray[87][242], dotarray[88][242], dotarray[89][242], dotarray[90][242], dotarray[91][242], dotarray[92][242], dotarray[93][242], dotarray[94][242], dotarray[95][242], dotarray[96][242], dotarray[97][242], dotarray[98][242], dotarray[99][242], dotarray[100][242], dotarray[101][242], dotarray[102][242], dotarray[103][242], dotarray[104][242], dotarray[105][242], dotarray[106][242], dotarray[107][242], dotarray[108][242], dotarray[109][242], dotarray[110][242], dotarray[111][242], dotarray[112][242], dotarray[113][242], dotarray[114][242], dotarray[115][242], dotarray[116][242], dotarray[117][242], dotarray[118][242], dotarray[119][242], dotarray[120][242], dotarray[121][242], dotarray[122][242], dotarray[123][242], dotarray[124][242], dotarray[125][242], dotarray[126][242], dotarray[127][242]};
assign dot_col_243 = {dotarray[0][243], dotarray[1][243], dotarray[2][243], dotarray[3][243], dotarray[4][243], dotarray[5][243], dotarray[6][243], dotarray[7][243], dotarray[8][243], dotarray[9][243], dotarray[10][243], dotarray[11][243], dotarray[12][243], dotarray[13][243], dotarray[14][243], dotarray[15][243], dotarray[16][243], dotarray[17][243], dotarray[18][243], dotarray[19][243], dotarray[20][243], dotarray[21][243], dotarray[22][243], dotarray[23][243], dotarray[24][243], dotarray[25][243], dotarray[26][243], dotarray[27][243], dotarray[28][243], dotarray[29][243], dotarray[30][243], dotarray[31][243], dotarray[32][243], dotarray[33][243], dotarray[34][243], dotarray[35][243], dotarray[36][243], dotarray[37][243], dotarray[38][243], dotarray[39][243], dotarray[40][243], dotarray[41][243], dotarray[42][243], dotarray[43][243], dotarray[44][243], dotarray[45][243], dotarray[46][243], dotarray[47][243], dotarray[48][243], dotarray[49][243], dotarray[50][243], dotarray[51][243], dotarray[52][243], dotarray[53][243], dotarray[54][243], dotarray[55][243], dotarray[56][243], dotarray[57][243], dotarray[58][243], dotarray[59][243], dotarray[60][243], dotarray[61][243], dotarray[62][243], dotarray[63][243], dotarray[64][243], dotarray[65][243], dotarray[66][243], dotarray[67][243], dotarray[68][243], dotarray[69][243], dotarray[70][243], dotarray[71][243], dotarray[72][243], dotarray[73][243], dotarray[74][243], dotarray[75][243], dotarray[76][243], dotarray[77][243], dotarray[78][243], dotarray[79][243], dotarray[80][243], dotarray[81][243], dotarray[82][243], dotarray[83][243], dotarray[84][243], dotarray[85][243], dotarray[86][243], dotarray[87][243], dotarray[88][243], dotarray[89][243], dotarray[90][243], dotarray[91][243], dotarray[92][243], dotarray[93][243], dotarray[94][243], dotarray[95][243], dotarray[96][243], dotarray[97][243], dotarray[98][243], dotarray[99][243], dotarray[100][243], dotarray[101][243], dotarray[102][243], dotarray[103][243], dotarray[104][243], dotarray[105][243], dotarray[106][243], dotarray[107][243], dotarray[108][243], dotarray[109][243], dotarray[110][243], dotarray[111][243], dotarray[112][243], dotarray[113][243], dotarray[114][243], dotarray[115][243], dotarray[116][243], dotarray[117][243], dotarray[118][243], dotarray[119][243], dotarray[120][243], dotarray[121][243], dotarray[122][243], dotarray[123][243], dotarray[124][243], dotarray[125][243], dotarray[126][243], dotarray[127][243]};
assign dot_col_244 = {dotarray[0][244], dotarray[1][244], dotarray[2][244], dotarray[3][244], dotarray[4][244], dotarray[5][244], dotarray[6][244], dotarray[7][244], dotarray[8][244], dotarray[9][244], dotarray[10][244], dotarray[11][244], dotarray[12][244], dotarray[13][244], dotarray[14][244], dotarray[15][244], dotarray[16][244], dotarray[17][244], dotarray[18][244], dotarray[19][244], dotarray[20][244], dotarray[21][244], dotarray[22][244], dotarray[23][244], dotarray[24][244], dotarray[25][244], dotarray[26][244], dotarray[27][244], dotarray[28][244], dotarray[29][244], dotarray[30][244], dotarray[31][244], dotarray[32][244], dotarray[33][244], dotarray[34][244], dotarray[35][244], dotarray[36][244], dotarray[37][244], dotarray[38][244], dotarray[39][244], dotarray[40][244], dotarray[41][244], dotarray[42][244], dotarray[43][244], dotarray[44][244], dotarray[45][244], dotarray[46][244], dotarray[47][244], dotarray[48][244], dotarray[49][244], dotarray[50][244], dotarray[51][244], dotarray[52][244], dotarray[53][244], dotarray[54][244], dotarray[55][244], dotarray[56][244], dotarray[57][244], dotarray[58][244], dotarray[59][244], dotarray[60][244], dotarray[61][244], dotarray[62][244], dotarray[63][244], dotarray[64][244], dotarray[65][244], dotarray[66][244], dotarray[67][244], dotarray[68][244], dotarray[69][244], dotarray[70][244], dotarray[71][244], dotarray[72][244], dotarray[73][244], dotarray[74][244], dotarray[75][244], dotarray[76][244], dotarray[77][244], dotarray[78][244], dotarray[79][244], dotarray[80][244], dotarray[81][244], dotarray[82][244], dotarray[83][244], dotarray[84][244], dotarray[85][244], dotarray[86][244], dotarray[87][244], dotarray[88][244], dotarray[89][244], dotarray[90][244], dotarray[91][244], dotarray[92][244], dotarray[93][244], dotarray[94][244], dotarray[95][244], dotarray[96][244], dotarray[97][244], dotarray[98][244], dotarray[99][244], dotarray[100][244], dotarray[101][244], dotarray[102][244], dotarray[103][244], dotarray[104][244], dotarray[105][244], dotarray[106][244], dotarray[107][244], dotarray[108][244], dotarray[109][244], dotarray[110][244], dotarray[111][244], dotarray[112][244], dotarray[113][244], dotarray[114][244], dotarray[115][244], dotarray[116][244], dotarray[117][244], dotarray[118][244], dotarray[119][244], dotarray[120][244], dotarray[121][244], dotarray[122][244], dotarray[123][244], dotarray[124][244], dotarray[125][244], dotarray[126][244], dotarray[127][244]};
assign dot_col_245 = {dotarray[0][245], dotarray[1][245], dotarray[2][245], dotarray[3][245], dotarray[4][245], dotarray[5][245], dotarray[6][245], dotarray[7][245], dotarray[8][245], dotarray[9][245], dotarray[10][245], dotarray[11][245], dotarray[12][245], dotarray[13][245], dotarray[14][245], dotarray[15][245], dotarray[16][245], dotarray[17][245], dotarray[18][245], dotarray[19][245], dotarray[20][245], dotarray[21][245], dotarray[22][245], dotarray[23][245], dotarray[24][245], dotarray[25][245], dotarray[26][245], dotarray[27][245], dotarray[28][245], dotarray[29][245], dotarray[30][245], dotarray[31][245], dotarray[32][245], dotarray[33][245], dotarray[34][245], dotarray[35][245], dotarray[36][245], dotarray[37][245], dotarray[38][245], dotarray[39][245], dotarray[40][245], dotarray[41][245], dotarray[42][245], dotarray[43][245], dotarray[44][245], dotarray[45][245], dotarray[46][245], dotarray[47][245], dotarray[48][245], dotarray[49][245], dotarray[50][245], dotarray[51][245], dotarray[52][245], dotarray[53][245], dotarray[54][245], dotarray[55][245], dotarray[56][245], dotarray[57][245], dotarray[58][245], dotarray[59][245], dotarray[60][245], dotarray[61][245], dotarray[62][245], dotarray[63][245], dotarray[64][245], dotarray[65][245], dotarray[66][245], dotarray[67][245], dotarray[68][245], dotarray[69][245], dotarray[70][245], dotarray[71][245], dotarray[72][245], dotarray[73][245], dotarray[74][245], dotarray[75][245], dotarray[76][245], dotarray[77][245], dotarray[78][245], dotarray[79][245], dotarray[80][245], dotarray[81][245], dotarray[82][245], dotarray[83][245], dotarray[84][245], dotarray[85][245], dotarray[86][245], dotarray[87][245], dotarray[88][245], dotarray[89][245], dotarray[90][245], dotarray[91][245], dotarray[92][245], dotarray[93][245], dotarray[94][245], dotarray[95][245], dotarray[96][245], dotarray[97][245], dotarray[98][245], dotarray[99][245], dotarray[100][245], dotarray[101][245], dotarray[102][245], dotarray[103][245], dotarray[104][245], dotarray[105][245], dotarray[106][245], dotarray[107][245], dotarray[108][245], dotarray[109][245], dotarray[110][245], dotarray[111][245], dotarray[112][245], dotarray[113][245], dotarray[114][245], dotarray[115][245], dotarray[116][245], dotarray[117][245], dotarray[118][245], dotarray[119][245], dotarray[120][245], dotarray[121][245], dotarray[122][245], dotarray[123][245], dotarray[124][245], dotarray[125][245], dotarray[126][245], dotarray[127][245]};
assign dot_col_246 = {dotarray[0][246], dotarray[1][246], dotarray[2][246], dotarray[3][246], dotarray[4][246], dotarray[5][246], dotarray[6][246], dotarray[7][246], dotarray[8][246], dotarray[9][246], dotarray[10][246], dotarray[11][246], dotarray[12][246], dotarray[13][246], dotarray[14][246], dotarray[15][246], dotarray[16][246], dotarray[17][246], dotarray[18][246], dotarray[19][246], dotarray[20][246], dotarray[21][246], dotarray[22][246], dotarray[23][246], dotarray[24][246], dotarray[25][246], dotarray[26][246], dotarray[27][246], dotarray[28][246], dotarray[29][246], dotarray[30][246], dotarray[31][246], dotarray[32][246], dotarray[33][246], dotarray[34][246], dotarray[35][246], dotarray[36][246], dotarray[37][246], dotarray[38][246], dotarray[39][246], dotarray[40][246], dotarray[41][246], dotarray[42][246], dotarray[43][246], dotarray[44][246], dotarray[45][246], dotarray[46][246], dotarray[47][246], dotarray[48][246], dotarray[49][246], dotarray[50][246], dotarray[51][246], dotarray[52][246], dotarray[53][246], dotarray[54][246], dotarray[55][246], dotarray[56][246], dotarray[57][246], dotarray[58][246], dotarray[59][246], dotarray[60][246], dotarray[61][246], dotarray[62][246], dotarray[63][246], dotarray[64][246], dotarray[65][246], dotarray[66][246], dotarray[67][246], dotarray[68][246], dotarray[69][246], dotarray[70][246], dotarray[71][246], dotarray[72][246], dotarray[73][246], dotarray[74][246], dotarray[75][246], dotarray[76][246], dotarray[77][246], dotarray[78][246], dotarray[79][246], dotarray[80][246], dotarray[81][246], dotarray[82][246], dotarray[83][246], dotarray[84][246], dotarray[85][246], dotarray[86][246], dotarray[87][246], dotarray[88][246], dotarray[89][246], dotarray[90][246], dotarray[91][246], dotarray[92][246], dotarray[93][246], dotarray[94][246], dotarray[95][246], dotarray[96][246], dotarray[97][246], dotarray[98][246], dotarray[99][246], dotarray[100][246], dotarray[101][246], dotarray[102][246], dotarray[103][246], dotarray[104][246], dotarray[105][246], dotarray[106][246], dotarray[107][246], dotarray[108][246], dotarray[109][246], dotarray[110][246], dotarray[111][246], dotarray[112][246], dotarray[113][246], dotarray[114][246], dotarray[115][246], dotarray[116][246], dotarray[117][246], dotarray[118][246], dotarray[119][246], dotarray[120][246], dotarray[121][246], dotarray[122][246], dotarray[123][246], dotarray[124][246], dotarray[125][246], dotarray[126][246], dotarray[127][246]};
assign dot_col_247 = {dotarray[0][247], dotarray[1][247], dotarray[2][247], dotarray[3][247], dotarray[4][247], dotarray[5][247], dotarray[6][247], dotarray[7][247], dotarray[8][247], dotarray[9][247], dotarray[10][247], dotarray[11][247], dotarray[12][247], dotarray[13][247], dotarray[14][247], dotarray[15][247], dotarray[16][247], dotarray[17][247], dotarray[18][247], dotarray[19][247], dotarray[20][247], dotarray[21][247], dotarray[22][247], dotarray[23][247], dotarray[24][247], dotarray[25][247], dotarray[26][247], dotarray[27][247], dotarray[28][247], dotarray[29][247], dotarray[30][247], dotarray[31][247], dotarray[32][247], dotarray[33][247], dotarray[34][247], dotarray[35][247], dotarray[36][247], dotarray[37][247], dotarray[38][247], dotarray[39][247], dotarray[40][247], dotarray[41][247], dotarray[42][247], dotarray[43][247], dotarray[44][247], dotarray[45][247], dotarray[46][247], dotarray[47][247], dotarray[48][247], dotarray[49][247], dotarray[50][247], dotarray[51][247], dotarray[52][247], dotarray[53][247], dotarray[54][247], dotarray[55][247], dotarray[56][247], dotarray[57][247], dotarray[58][247], dotarray[59][247], dotarray[60][247], dotarray[61][247], dotarray[62][247], dotarray[63][247], dotarray[64][247], dotarray[65][247], dotarray[66][247], dotarray[67][247], dotarray[68][247], dotarray[69][247], dotarray[70][247], dotarray[71][247], dotarray[72][247], dotarray[73][247], dotarray[74][247], dotarray[75][247], dotarray[76][247], dotarray[77][247], dotarray[78][247], dotarray[79][247], dotarray[80][247], dotarray[81][247], dotarray[82][247], dotarray[83][247], dotarray[84][247], dotarray[85][247], dotarray[86][247], dotarray[87][247], dotarray[88][247], dotarray[89][247], dotarray[90][247], dotarray[91][247], dotarray[92][247], dotarray[93][247], dotarray[94][247], dotarray[95][247], dotarray[96][247], dotarray[97][247], dotarray[98][247], dotarray[99][247], dotarray[100][247], dotarray[101][247], dotarray[102][247], dotarray[103][247], dotarray[104][247], dotarray[105][247], dotarray[106][247], dotarray[107][247], dotarray[108][247], dotarray[109][247], dotarray[110][247], dotarray[111][247], dotarray[112][247], dotarray[113][247], dotarray[114][247], dotarray[115][247], dotarray[116][247], dotarray[117][247], dotarray[118][247], dotarray[119][247], dotarray[120][247], dotarray[121][247], dotarray[122][247], dotarray[123][247], dotarray[124][247], dotarray[125][247], dotarray[126][247], dotarray[127][247]};
assign dot_col_248 = {dotarray[0][248], dotarray[1][248], dotarray[2][248], dotarray[3][248], dotarray[4][248], dotarray[5][248], dotarray[6][248], dotarray[7][248], dotarray[8][248], dotarray[9][248], dotarray[10][248], dotarray[11][248], dotarray[12][248], dotarray[13][248], dotarray[14][248], dotarray[15][248], dotarray[16][248], dotarray[17][248], dotarray[18][248], dotarray[19][248], dotarray[20][248], dotarray[21][248], dotarray[22][248], dotarray[23][248], dotarray[24][248], dotarray[25][248], dotarray[26][248], dotarray[27][248], dotarray[28][248], dotarray[29][248], dotarray[30][248], dotarray[31][248], dotarray[32][248], dotarray[33][248], dotarray[34][248], dotarray[35][248], dotarray[36][248], dotarray[37][248], dotarray[38][248], dotarray[39][248], dotarray[40][248], dotarray[41][248], dotarray[42][248], dotarray[43][248], dotarray[44][248], dotarray[45][248], dotarray[46][248], dotarray[47][248], dotarray[48][248], dotarray[49][248], dotarray[50][248], dotarray[51][248], dotarray[52][248], dotarray[53][248], dotarray[54][248], dotarray[55][248], dotarray[56][248], dotarray[57][248], dotarray[58][248], dotarray[59][248], dotarray[60][248], dotarray[61][248], dotarray[62][248], dotarray[63][248], dotarray[64][248], dotarray[65][248], dotarray[66][248], dotarray[67][248], dotarray[68][248], dotarray[69][248], dotarray[70][248], dotarray[71][248], dotarray[72][248], dotarray[73][248], dotarray[74][248], dotarray[75][248], dotarray[76][248], dotarray[77][248], dotarray[78][248], dotarray[79][248], dotarray[80][248], dotarray[81][248], dotarray[82][248], dotarray[83][248], dotarray[84][248], dotarray[85][248], dotarray[86][248], dotarray[87][248], dotarray[88][248], dotarray[89][248], dotarray[90][248], dotarray[91][248], dotarray[92][248], dotarray[93][248], dotarray[94][248], dotarray[95][248], dotarray[96][248], dotarray[97][248], dotarray[98][248], dotarray[99][248], dotarray[100][248], dotarray[101][248], dotarray[102][248], dotarray[103][248], dotarray[104][248], dotarray[105][248], dotarray[106][248], dotarray[107][248], dotarray[108][248], dotarray[109][248], dotarray[110][248], dotarray[111][248], dotarray[112][248], dotarray[113][248], dotarray[114][248], dotarray[115][248], dotarray[116][248], dotarray[117][248], dotarray[118][248], dotarray[119][248], dotarray[120][248], dotarray[121][248], dotarray[122][248], dotarray[123][248], dotarray[124][248], dotarray[125][248], dotarray[126][248], dotarray[127][248]};
assign dot_col_249 = {dotarray[0][249], dotarray[1][249], dotarray[2][249], dotarray[3][249], dotarray[4][249], dotarray[5][249], dotarray[6][249], dotarray[7][249], dotarray[8][249], dotarray[9][249], dotarray[10][249], dotarray[11][249], dotarray[12][249], dotarray[13][249], dotarray[14][249], dotarray[15][249], dotarray[16][249], dotarray[17][249], dotarray[18][249], dotarray[19][249], dotarray[20][249], dotarray[21][249], dotarray[22][249], dotarray[23][249], dotarray[24][249], dotarray[25][249], dotarray[26][249], dotarray[27][249], dotarray[28][249], dotarray[29][249], dotarray[30][249], dotarray[31][249], dotarray[32][249], dotarray[33][249], dotarray[34][249], dotarray[35][249], dotarray[36][249], dotarray[37][249], dotarray[38][249], dotarray[39][249], dotarray[40][249], dotarray[41][249], dotarray[42][249], dotarray[43][249], dotarray[44][249], dotarray[45][249], dotarray[46][249], dotarray[47][249], dotarray[48][249], dotarray[49][249], dotarray[50][249], dotarray[51][249], dotarray[52][249], dotarray[53][249], dotarray[54][249], dotarray[55][249], dotarray[56][249], dotarray[57][249], dotarray[58][249], dotarray[59][249], dotarray[60][249], dotarray[61][249], dotarray[62][249], dotarray[63][249], dotarray[64][249], dotarray[65][249], dotarray[66][249], dotarray[67][249], dotarray[68][249], dotarray[69][249], dotarray[70][249], dotarray[71][249], dotarray[72][249], dotarray[73][249], dotarray[74][249], dotarray[75][249], dotarray[76][249], dotarray[77][249], dotarray[78][249], dotarray[79][249], dotarray[80][249], dotarray[81][249], dotarray[82][249], dotarray[83][249], dotarray[84][249], dotarray[85][249], dotarray[86][249], dotarray[87][249], dotarray[88][249], dotarray[89][249], dotarray[90][249], dotarray[91][249], dotarray[92][249], dotarray[93][249], dotarray[94][249], dotarray[95][249], dotarray[96][249], dotarray[97][249], dotarray[98][249], dotarray[99][249], dotarray[100][249], dotarray[101][249], dotarray[102][249], dotarray[103][249], dotarray[104][249], dotarray[105][249], dotarray[106][249], dotarray[107][249], dotarray[108][249], dotarray[109][249], dotarray[110][249], dotarray[111][249], dotarray[112][249], dotarray[113][249], dotarray[114][249], dotarray[115][249], dotarray[116][249], dotarray[117][249], dotarray[118][249], dotarray[119][249], dotarray[120][249], dotarray[121][249], dotarray[122][249], dotarray[123][249], dotarray[124][249], dotarray[125][249], dotarray[126][249], dotarray[127][249]};
assign dot_col_250 = {dotarray[0][250], dotarray[1][250], dotarray[2][250], dotarray[3][250], dotarray[4][250], dotarray[5][250], dotarray[6][250], dotarray[7][250], dotarray[8][250], dotarray[9][250], dotarray[10][250], dotarray[11][250], dotarray[12][250], dotarray[13][250], dotarray[14][250], dotarray[15][250], dotarray[16][250], dotarray[17][250], dotarray[18][250], dotarray[19][250], dotarray[20][250], dotarray[21][250], dotarray[22][250], dotarray[23][250], dotarray[24][250], dotarray[25][250], dotarray[26][250], dotarray[27][250], dotarray[28][250], dotarray[29][250], dotarray[30][250], dotarray[31][250], dotarray[32][250], dotarray[33][250], dotarray[34][250], dotarray[35][250], dotarray[36][250], dotarray[37][250], dotarray[38][250], dotarray[39][250], dotarray[40][250], dotarray[41][250], dotarray[42][250], dotarray[43][250], dotarray[44][250], dotarray[45][250], dotarray[46][250], dotarray[47][250], dotarray[48][250], dotarray[49][250], dotarray[50][250], dotarray[51][250], dotarray[52][250], dotarray[53][250], dotarray[54][250], dotarray[55][250], dotarray[56][250], dotarray[57][250], dotarray[58][250], dotarray[59][250], dotarray[60][250], dotarray[61][250], dotarray[62][250], dotarray[63][250], dotarray[64][250], dotarray[65][250], dotarray[66][250], dotarray[67][250], dotarray[68][250], dotarray[69][250], dotarray[70][250], dotarray[71][250], dotarray[72][250], dotarray[73][250], dotarray[74][250], dotarray[75][250], dotarray[76][250], dotarray[77][250], dotarray[78][250], dotarray[79][250], dotarray[80][250], dotarray[81][250], dotarray[82][250], dotarray[83][250], dotarray[84][250], dotarray[85][250], dotarray[86][250], dotarray[87][250], dotarray[88][250], dotarray[89][250], dotarray[90][250], dotarray[91][250], dotarray[92][250], dotarray[93][250], dotarray[94][250], dotarray[95][250], dotarray[96][250], dotarray[97][250], dotarray[98][250], dotarray[99][250], dotarray[100][250], dotarray[101][250], dotarray[102][250], dotarray[103][250], dotarray[104][250], dotarray[105][250], dotarray[106][250], dotarray[107][250], dotarray[108][250], dotarray[109][250], dotarray[110][250], dotarray[111][250], dotarray[112][250], dotarray[113][250], dotarray[114][250], dotarray[115][250], dotarray[116][250], dotarray[117][250], dotarray[118][250], dotarray[119][250], dotarray[120][250], dotarray[121][250], dotarray[122][250], dotarray[123][250], dotarray[124][250], dotarray[125][250], dotarray[126][250], dotarray[127][250]};
assign dot_col_251 = {dotarray[0][251], dotarray[1][251], dotarray[2][251], dotarray[3][251], dotarray[4][251], dotarray[5][251], dotarray[6][251], dotarray[7][251], dotarray[8][251], dotarray[9][251], dotarray[10][251], dotarray[11][251], dotarray[12][251], dotarray[13][251], dotarray[14][251], dotarray[15][251], dotarray[16][251], dotarray[17][251], dotarray[18][251], dotarray[19][251], dotarray[20][251], dotarray[21][251], dotarray[22][251], dotarray[23][251], dotarray[24][251], dotarray[25][251], dotarray[26][251], dotarray[27][251], dotarray[28][251], dotarray[29][251], dotarray[30][251], dotarray[31][251], dotarray[32][251], dotarray[33][251], dotarray[34][251], dotarray[35][251], dotarray[36][251], dotarray[37][251], dotarray[38][251], dotarray[39][251], dotarray[40][251], dotarray[41][251], dotarray[42][251], dotarray[43][251], dotarray[44][251], dotarray[45][251], dotarray[46][251], dotarray[47][251], dotarray[48][251], dotarray[49][251], dotarray[50][251], dotarray[51][251], dotarray[52][251], dotarray[53][251], dotarray[54][251], dotarray[55][251], dotarray[56][251], dotarray[57][251], dotarray[58][251], dotarray[59][251], dotarray[60][251], dotarray[61][251], dotarray[62][251], dotarray[63][251], dotarray[64][251], dotarray[65][251], dotarray[66][251], dotarray[67][251], dotarray[68][251], dotarray[69][251], dotarray[70][251], dotarray[71][251], dotarray[72][251], dotarray[73][251], dotarray[74][251], dotarray[75][251], dotarray[76][251], dotarray[77][251], dotarray[78][251], dotarray[79][251], dotarray[80][251], dotarray[81][251], dotarray[82][251], dotarray[83][251], dotarray[84][251], dotarray[85][251], dotarray[86][251], dotarray[87][251], dotarray[88][251], dotarray[89][251], dotarray[90][251], dotarray[91][251], dotarray[92][251], dotarray[93][251], dotarray[94][251], dotarray[95][251], dotarray[96][251], dotarray[97][251], dotarray[98][251], dotarray[99][251], dotarray[100][251], dotarray[101][251], dotarray[102][251], dotarray[103][251], dotarray[104][251], dotarray[105][251], dotarray[106][251], dotarray[107][251], dotarray[108][251], dotarray[109][251], dotarray[110][251], dotarray[111][251], dotarray[112][251], dotarray[113][251], dotarray[114][251], dotarray[115][251], dotarray[116][251], dotarray[117][251], dotarray[118][251], dotarray[119][251], dotarray[120][251], dotarray[121][251], dotarray[122][251], dotarray[123][251], dotarray[124][251], dotarray[125][251], dotarray[126][251], dotarray[127][251]};
assign dot_col_252 = {dotarray[0][252], dotarray[1][252], dotarray[2][252], dotarray[3][252], dotarray[4][252], dotarray[5][252], dotarray[6][252], dotarray[7][252], dotarray[8][252], dotarray[9][252], dotarray[10][252], dotarray[11][252], dotarray[12][252], dotarray[13][252], dotarray[14][252], dotarray[15][252], dotarray[16][252], dotarray[17][252], dotarray[18][252], dotarray[19][252], dotarray[20][252], dotarray[21][252], dotarray[22][252], dotarray[23][252], dotarray[24][252], dotarray[25][252], dotarray[26][252], dotarray[27][252], dotarray[28][252], dotarray[29][252], dotarray[30][252], dotarray[31][252], dotarray[32][252], dotarray[33][252], dotarray[34][252], dotarray[35][252], dotarray[36][252], dotarray[37][252], dotarray[38][252], dotarray[39][252], dotarray[40][252], dotarray[41][252], dotarray[42][252], dotarray[43][252], dotarray[44][252], dotarray[45][252], dotarray[46][252], dotarray[47][252], dotarray[48][252], dotarray[49][252], dotarray[50][252], dotarray[51][252], dotarray[52][252], dotarray[53][252], dotarray[54][252], dotarray[55][252], dotarray[56][252], dotarray[57][252], dotarray[58][252], dotarray[59][252], dotarray[60][252], dotarray[61][252], dotarray[62][252], dotarray[63][252], dotarray[64][252], dotarray[65][252], dotarray[66][252], dotarray[67][252], dotarray[68][252], dotarray[69][252], dotarray[70][252], dotarray[71][252], dotarray[72][252], dotarray[73][252], dotarray[74][252], dotarray[75][252], dotarray[76][252], dotarray[77][252], dotarray[78][252], dotarray[79][252], dotarray[80][252], dotarray[81][252], dotarray[82][252], dotarray[83][252], dotarray[84][252], dotarray[85][252], dotarray[86][252], dotarray[87][252], dotarray[88][252], dotarray[89][252], dotarray[90][252], dotarray[91][252], dotarray[92][252], dotarray[93][252], dotarray[94][252], dotarray[95][252], dotarray[96][252], dotarray[97][252], dotarray[98][252], dotarray[99][252], dotarray[100][252], dotarray[101][252], dotarray[102][252], dotarray[103][252], dotarray[104][252], dotarray[105][252], dotarray[106][252], dotarray[107][252], dotarray[108][252], dotarray[109][252], dotarray[110][252], dotarray[111][252], dotarray[112][252], dotarray[113][252], dotarray[114][252], dotarray[115][252], dotarray[116][252], dotarray[117][252], dotarray[118][252], dotarray[119][252], dotarray[120][252], dotarray[121][252], dotarray[122][252], dotarray[123][252], dotarray[124][252], dotarray[125][252], dotarray[126][252], dotarray[127][252]};
assign dot_col_253 = {dotarray[0][253], dotarray[1][253], dotarray[2][253], dotarray[3][253], dotarray[4][253], dotarray[5][253], dotarray[6][253], dotarray[7][253], dotarray[8][253], dotarray[9][253], dotarray[10][253], dotarray[11][253], dotarray[12][253], dotarray[13][253], dotarray[14][253], dotarray[15][253], dotarray[16][253], dotarray[17][253], dotarray[18][253], dotarray[19][253], dotarray[20][253], dotarray[21][253], dotarray[22][253], dotarray[23][253], dotarray[24][253], dotarray[25][253], dotarray[26][253], dotarray[27][253], dotarray[28][253], dotarray[29][253], dotarray[30][253], dotarray[31][253], dotarray[32][253], dotarray[33][253], dotarray[34][253], dotarray[35][253], dotarray[36][253], dotarray[37][253], dotarray[38][253], dotarray[39][253], dotarray[40][253], dotarray[41][253], dotarray[42][253], dotarray[43][253], dotarray[44][253], dotarray[45][253], dotarray[46][253], dotarray[47][253], dotarray[48][253], dotarray[49][253], dotarray[50][253], dotarray[51][253], dotarray[52][253], dotarray[53][253], dotarray[54][253], dotarray[55][253], dotarray[56][253], dotarray[57][253], dotarray[58][253], dotarray[59][253], dotarray[60][253], dotarray[61][253], dotarray[62][253], dotarray[63][253], dotarray[64][253], dotarray[65][253], dotarray[66][253], dotarray[67][253], dotarray[68][253], dotarray[69][253], dotarray[70][253], dotarray[71][253], dotarray[72][253], dotarray[73][253], dotarray[74][253], dotarray[75][253], dotarray[76][253], dotarray[77][253], dotarray[78][253], dotarray[79][253], dotarray[80][253], dotarray[81][253], dotarray[82][253], dotarray[83][253], dotarray[84][253], dotarray[85][253], dotarray[86][253], dotarray[87][253], dotarray[88][253], dotarray[89][253], dotarray[90][253], dotarray[91][253], dotarray[92][253], dotarray[93][253], dotarray[94][253], dotarray[95][253], dotarray[96][253], dotarray[97][253], dotarray[98][253], dotarray[99][253], dotarray[100][253], dotarray[101][253], dotarray[102][253], dotarray[103][253], dotarray[104][253], dotarray[105][253], dotarray[106][253], dotarray[107][253], dotarray[108][253], dotarray[109][253], dotarray[110][253], dotarray[111][253], dotarray[112][253], dotarray[113][253], dotarray[114][253], dotarray[115][253], dotarray[116][253], dotarray[117][253], dotarray[118][253], dotarray[119][253], dotarray[120][253], dotarray[121][253], dotarray[122][253], dotarray[123][253], dotarray[124][253], dotarray[125][253], dotarray[126][253], dotarray[127][253]};
assign dot_col_254 = {dotarray[0][254], dotarray[1][254], dotarray[2][254], dotarray[3][254], dotarray[4][254], dotarray[5][254], dotarray[6][254], dotarray[7][254], dotarray[8][254], dotarray[9][254], dotarray[10][254], dotarray[11][254], dotarray[12][254], dotarray[13][254], dotarray[14][254], dotarray[15][254], dotarray[16][254], dotarray[17][254], dotarray[18][254], dotarray[19][254], dotarray[20][254], dotarray[21][254], dotarray[22][254], dotarray[23][254], dotarray[24][254], dotarray[25][254], dotarray[26][254], dotarray[27][254], dotarray[28][254], dotarray[29][254], dotarray[30][254], dotarray[31][254], dotarray[32][254], dotarray[33][254], dotarray[34][254], dotarray[35][254], dotarray[36][254], dotarray[37][254], dotarray[38][254], dotarray[39][254], dotarray[40][254], dotarray[41][254], dotarray[42][254], dotarray[43][254], dotarray[44][254], dotarray[45][254], dotarray[46][254], dotarray[47][254], dotarray[48][254], dotarray[49][254], dotarray[50][254], dotarray[51][254], dotarray[52][254], dotarray[53][254], dotarray[54][254], dotarray[55][254], dotarray[56][254], dotarray[57][254], dotarray[58][254], dotarray[59][254], dotarray[60][254], dotarray[61][254], dotarray[62][254], dotarray[63][254], dotarray[64][254], dotarray[65][254], dotarray[66][254], dotarray[67][254], dotarray[68][254], dotarray[69][254], dotarray[70][254], dotarray[71][254], dotarray[72][254], dotarray[73][254], dotarray[74][254], dotarray[75][254], dotarray[76][254], dotarray[77][254], dotarray[78][254], dotarray[79][254], dotarray[80][254], dotarray[81][254], dotarray[82][254], dotarray[83][254], dotarray[84][254], dotarray[85][254], dotarray[86][254], dotarray[87][254], dotarray[88][254], dotarray[89][254], dotarray[90][254], dotarray[91][254], dotarray[92][254], dotarray[93][254], dotarray[94][254], dotarray[95][254], dotarray[96][254], dotarray[97][254], dotarray[98][254], dotarray[99][254], dotarray[100][254], dotarray[101][254], dotarray[102][254], dotarray[103][254], dotarray[104][254], dotarray[105][254], dotarray[106][254], dotarray[107][254], dotarray[108][254], dotarray[109][254], dotarray[110][254], dotarray[111][254], dotarray[112][254], dotarray[113][254], dotarray[114][254], dotarray[115][254], dotarray[116][254], dotarray[117][254], dotarray[118][254], dotarray[119][254], dotarray[120][254], dotarray[121][254], dotarray[122][254], dotarray[123][254], dotarray[124][254], dotarray[125][254], dotarray[126][254], dotarray[127][254]};
assign dot_col_255 = {dotarray[0][255], dotarray[1][255], dotarray[2][255], dotarray[3][255], dotarray[4][255], dotarray[5][255], dotarray[6][255], dotarray[7][255], dotarray[8][255], dotarray[9][255], dotarray[10][255], dotarray[11][255], dotarray[12][255], dotarray[13][255], dotarray[14][255], dotarray[15][255], dotarray[16][255], dotarray[17][255], dotarray[18][255], dotarray[19][255], dotarray[20][255], dotarray[21][255], dotarray[22][255], dotarray[23][255], dotarray[24][255], dotarray[25][255], dotarray[26][255], dotarray[27][255], dotarray[28][255], dotarray[29][255], dotarray[30][255], dotarray[31][255], dotarray[32][255], dotarray[33][255], dotarray[34][255], dotarray[35][255], dotarray[36][255], dotarray[37][255], dotarray[38][255], dotarray[39][255], dotarray[40][255], dotarray[41][255], dotarray[42][255], dotarray[43][255], dotarray[44][255], dotarray[45][255], dotarray[46][255], dotarray[47][255], dotarray[48][255], dotarray[49][255], dotarray[50][255], dotarray[51][255], dotarray[52][255], dotarray[53][255], dotarray[54][255], dotarray[55][255], dotarray[56][255], dotarray[57][255], dotarray[58][255], dotarray[59][255], dotarray[60][255], dotarray[61][255], dotarray[62][255], dotarray[63][255], dotarray[64][255], dotarray[65][255], dotarray[66][255], dotarray[67][255], dotarray[68][255], dotarray[69][255], dotarray[70][255], dotarray[71][255], dotarray[72][255], dotarray[73][255], dotarray[74][255], dotarray[75][255], dotarray[76][255], dotarray[77][255], dotarray[78][255], dotarray[79][255], dotarray[80][255], dotarray[81][255], dotarray[82][255], dotarray[83][255], dotarray[84][255], dotarray[85][255], dotarray[86][255], dotarray[87][255], dotarray[88][255], dotarray[89][255], dotarray[90][255], dotarray[91][255], dotarray[92][255], dotarray[93][255], dotarray[94][255], dotarray[95][255], dotarray[96][255], dotarray[97][255], dotarray[98][255], dotarray[99][255], dotarray[100][255], dotarray[101][255], dotarray[102][255], dotarray[103][255], dotarray[104][255], dotarray[105][255], dotarray[106][255], dotarray[107][255], dotarray[108][255], dotarray[109][255], dotarray[110][255], dotarray[111][255], dotarray[112][255], dotarray[113][255], dotarray[114][255], dotarray[115][255], dotarray[116][255], dotarray[117][255], dotarray[118][255], dotarray[119][255], dotarray[120][255], dotarray[121][255], dotarray[122][255], dotarray[123][255], dotarray[124][255], dotarray[125][255], dotarray[126][255], dotarray[127][255]};

wire [7:0] check_col_0, check_col_1, check_col_2, check_col_3, check_col_4, check_col_5, check_col_6, check_col_7, 
           check_col_8, check_col_9, check_col_10, check_col_11, check_col_12, check_col_13, check_col_14, check_col_15, 
           check_col_16, check_col_17, check_col_18, check_col_19, check_col_20, check_col_21, check_col_22, check_col_23, 
           check_col_24, check_col_25, check_col_26, check_col_27, check_col_28, check_col_29, check_col_30, check_col_31, 
           check_col_32, check_col_33, check_col_34, check_col_35, check_col_36, check_col_37, check_col_38, check_col_39, 
           check_col_40, check_col_41, check_col_42, check_col_43, check_col_44, check_col_45, check_col_46, check_col_47, 
           check_col_48, check_col_49, check_col_50, check_col_51, check_col_52, check_col_53, check_col_54, check_col_55, 
           check_col_56, check_col_57, check_col_58, check_col_59, check_col_60, check_col_61, check_col_62, check_col_63, 
           check_col_64, check_col_65, check_col_66, check_col_67, check_col_68, check_col_69, check_col_70, check_col_71, 
           check_col_72, check_col_73, check_col_74, check_col_75, check_col_76, check_col_77, check_col_78, check_col_79, 
           check_col_80, check_col_81, check_col_82, check_col_83, check_col_84, check_col_85, check_col_86, check_col_87, 
           check_col_88, check_col_89, check_col_90, check_col_91, check_col_92, check_col_93, check_col_94, check_col_95, 
           check_col_96, check_col_97, check_col_98, check_col_99, check_col_100, check_col_101, check_col_102, check_col_103, 
           check_col_104, check_col_105, check_col_106, check_col_107, check_col_108, check_col_109, check_col_110, check_col_111, 
           check_col_112, check_col_113, check_col_114, check_col_115, check_col_116, check_col_117, check_col_118, check_col_119, 
           check_col_120, check_col_121, check_col_122, check_col_123, check_col_124, check_col_125, check_col_126, check_col_127, 
           check_col_128, check_col_129, check_col_130, check_col_131, check_col_132, check_col_133, check_col_134, check_col_135, 
           check_col_136, check_col_137, check_col_138, check_col_139, check_col_140, check_col_141, check_col_142, check_col_143, 
           check_col_144, check_col_145, check_col_146, check_col_147, check_col_148, check_col_149, check_col_150, check_col_151, 
           check_col_152, check_col_153, check_col_154, check_col_155, check_col_156, check_col_157, check_col_158, check_col_159, 
           check_col_160, check_col_161, check_col_162, check_col_163, check_col_164, check_col_165, check_col_166, check_col_167, 
           check_col_168, check_col_169, check_col_170, check_col_171, check_col_172, check_col_173, check_col_174, check_col_175, 
           check_col_176, check_col_177, check_col_178, check_col_179, check_col_180, check_col_181, check_col_182, check_col_183, 
           check_col_184, check_col_185, check_col_186, check_col_187, check_col_188, check_col_189, check_col_190, check_col_191, 
           check_col_192, check_col_193, check_col_194, check_col_195, check_col_196, check_col_197, check_col_198, check_col_199, 
           check_col_200, check_col_201, check_col_202, check_col_203, check_col_204, check_col_205, check_col_206, check_col_207, 
           check_col_208, check_col_209, check_col_210, check_col_211, check_col_212, check_col_213, check_col_214, check_col_215, 
           check_col_216, check_col_217, check_col_218, check_col_219, check_col_220, check_col_221, check_col_222, check_col_223, 
           check_col_224, check_col_225, check_col_226, check_col_227, check_col_228, check_col_229, check_col_230, check_col_231, 
           check_col_232, check_col_233, check_col_234, check_col_235, check_col_236, check_col_237, check_col_238, check_col_239, 
           check_col_240, check_col_241, check_col_242, check_col_243, check_col_244, check_col_245, check_col_246, check_col_247, 
           check_col_248, check_col_249, check_col_250, check_col_251, check_col_252, check_col_253, check_col_254, check_col_255;

wire [7:0] wrong_col_0, wrong_col_1, wrong_col_2, wrong_col_3, wrong_col_4, wrong_col_5, wrong_col_6, wrong_col_7, 
           wrong_col_8, wrong_col_9, wrong_col_10, wrong_col_11, wrong_col_12, wrong_col_13, wrong_col_14, wrong_col_15, 
           wrong_col_16, wrong_col_17, wrong_col_18, wrong_col_19, wrong_col_20, wrong_col_21, wrong_col_22, wrong_col_23, 
           wrong_col_24, wrong_col_25, wrong_col_26, wrong_col_27, wrong_col_28, wrong_col_29, wrong_col_30, wrong_col_31, 
           wrong_col_32, wrong_col_33, wrong_col_34, wrong_col_35, wrong_col_36, wrong_col_37, wrong_col_38, wrong_col_39, 
           wrong_col_40, wrong_col_41, wrong_col_42, wrong_col_43, wrong_col_44, wrong_col_45, wrong_col_46, wrong_col_47, 
           wrong_col_48, wrong_col_49, wrong_col_50, wrong_col_51, wrong_col_52, wrong_col_53, wrong_col_54, wrong_col_55, 
           wrong_col_56, wrong_col_57, wrong_col_58, wrong_col_59, wrong_col_60, wrong_col_61, wrong_col_62, wrong_col_63, 
           wrong_col_64, wrong_col_65, wrong_col_66, wrong_col_67, wrong_col_68, wrong_col_69, wrong_col_70, wrong_col_71, 
           wrong_col_72, wrong_col_73, wrong_col_74, wrong_col_75, wrong_col_76, wrong_col_77, wrong_col_78, wrong_col_79, 
           wrong_col_80, wrong_col_81, wrong_col_82, wrong_col_83, wrong_col_84, wrong_col_85, wrong_col_86, wrong_col_87, 
           wrong_col_88, wrong_col_89, wrong_col_90, wrong_col_91, wrong_col_92, wrong_col_93, wrong_col_94, wrong_col_95, 
           wrong_col_96, wrong_col_97, wrong_col_98, wrong_col_99, wrong_col_100, wrong_col_101, wrong_col_102, wrong_col_103, 
           wrong_col_104, wrong_col_105, wrong_col_106, wrong_col_107, wrong_col_108, wrong_col_109, wrong_col_110, wrong_col_111, 
           wrong_col_112, wrong_col_113, wrong_col_114, wrong_col_115, wrong_col_116, wrong_col_117, wrong_col_118, wrong_col_119, 
           wrong_col_120, wrong_col_121, wrong_col_122, wrong_col_123, wrong_col_124, wrong_col_125, wrong_col_126, wrong_col_127, 
           wrong_col_128, wrong_col_129, wrong_col_130, wrong_col_131, wrong_col_132, wrong_col_133, wrong_col_134, wrong_col_135, 
           wrong_col_136, wrong_col_137, wrong_col_138, wrong_col_139, wrong_col_140, wrong_col_141, wrong_col_142, wrong_col_143, 
           wrong_col_144, wrong_col_145, wrong_col_146, wrong_col_147, wrong_col_148, wrong_col_149, wrong_col_150, wrong_col_151, 
           wrong_col_152, wrong_col_153, wrong_col_154, wrong_col_155, wrong_col_156, wrong_col_157, wrong_col_158, wrong_col_159, 
           wrong_col_160, wrong_col_161, wrong_col_162, wrong_col_163, wrong_col_164, wrong_col_165, wrong_col_166, wrong_col_167, 
           wrong_col_168, wrong_col_169, wrong_col_170, wrong_col_171, wrong_col_172, wrong_col_173, wrong_col_174, wrong_col_175, 
           wrong_col_176, wrong_col_177, wrong_col_178, wrong_col_179, wrong_col_180, wrong_col_181, wrong_col_182, wrong_col_183, 
           wrong_col_184, wrong_col_185, wrong_col_186, wrong_col_187, wrong_col_188, wrong_col_189, wrong_col_190, wrong_col_191, 
           wrong_col_192, wrong_col_193, wrong_col_194, wrong_col_195, wrong_col_196, wrong_col_197, wrong_col_198, wrong_col_199, 
           wrong_col_200, wrong_col_201, wrong_col_202, wrong_col_203, wrong_col_204, wrong_col_205, wrong_col_206, wrong_col_207, 
           wrong_col_208, wrong_col_209, wrong_col_210, wrong_col_211, wrong_col_212, wrong_col_213, wrong_col_214, wrong_col_215, 
           wrong_col_216, wrong_col_217, wrong_col_218, wrong_col_219, wrong_col_220, wrong_col_221, wrong_col_222, wrong_col_223, 
           wrong_col_224, wrong_col_225, wrong_col_226, wrong_col_227, wrong_col_228, wrong_col_229, wrong_col_230, wrong_col_231, 
           wrong_col_232, wrong_col_233, wrong_col_234, wrong_col_235, wrong_col_236, wrong_col_237, wrong_col_238, wrong_col_239, 
           wrong_col_240, wrong_col_241, wrong_col_242, wrong_col_243, wrong_col_244, wrong_col_245, wrong_col_246, wrong_col_247, 
           wrong_col_248, wrong_col_249, wrong_col_250, wrong_col_251, wrong_col_252, wrong_col_253, wrong_col_254, wrong_col_255;

bitsadder_128 c_num_0(.data_in(dot_col_0), .sum(check_col_0));
bitsadder_128 c_num_1(.data_in(dot_col_1), .sum(check_col_1));
bitsadder_128 c_num_2(.data_in(dot_col_2), .sum(check_col_2));
bitsadder_128 c_num_3(.data_in(dot_col_3), .sum(check_col_3));
bitsadder_128 c_num_4(.data_in(dot_col_4), .sum(check_col_4));
bitsadder_128 c_num_5(.data_in(dot_col_5), .sum(check_col_5));
bitsadder_128 c_num_6(.data_in(dot_col_6), .sum(check_col_6));
bitsadder_128 c_num_7(.data_in(dot_col_7), .sum(check_col_7));
bitsadder_128 c_num_8(.data_in(dot_col_8), .sum(check_col_8));
bitsadder_128 c_num_9(.data_in(dot_col_9), .sum(check_col_9));
bitsadder_128 c_num_10(.data_in(dot_col_10), .sum(check_col_10));
bitsadder_128 c_num_11(.data_in(dot_col_11), .sum(check_col_11));
bitsadder_128 c_num_12(.data_in(dot_col_12), .sum(check_col_12));
bitsadder_128 c_num_13(.data_in(dot_col_13), .sum(check_col_13));
bitsadder_128 c_num_14(.data_in(dot_col_14), .sum(check_col_14));
bitsadder_128 c_num_15(.data_in(dot_col_15), .sum(check_col_15));
bitsadder_128 c_num_16(.data_in(dot_col_16), .sum(check_col_16));
bitsadder_128 c_num_17(.data_in(dot_col_17), .sum(check_col_17));
bitsadder_128 c_num_18(.data_in(dot_col_18), .sum(check_col_18));
bitsadder_128 c_num_19(.data_in(dot_col_19), .sum(check_col_19));
bitsadder_128 c_num_20(.data_in(dot_col_20), .sum(check_col_20));
bitsadder_128 c_num_21(.data_in(dot_col_21), .sum(check_col_21));
bitsadder_128 c_num_22(.data_in(dot_col_22), .sum(check_col_22));
bitsadder_128 c_num_23(.data_in(dot_col_23), .sum(check_col_23));
bitsadder_128 c_num_24(.data_in(dot_col_24), .sum(check_col_24));
bitsadder_128 c_num_25(.data_in(dot_col_25), .sum(check_col_25));
bitsadder_128 c_num_26(.data_in(dot_col_26), .sum(check_col_26));
bitsadder_128 c_num_27(.data_in(dot_col_27), .sum(check_col_27));
bitsadder_128 c_num_28(.data_in(dot_col_28), .sum(check_col_28));
bitsadder_128 c_num_29(.data_in(dot_col_29), .sum(check_col_29));
bitsadder_128 c_num_30(.data_in(dot_col_30), .sum(check_col_30));
bitsadder_128 c_num_31(.data_in(dot_col_31), .sum(check_col_31));
bitsadder_128 c_num_32(.data_in(dot_col_32), .sum(check_col_32));
bitsadder_128 c_num_33(.data_in(dot_col_33), .sum(check_col_33));
bitsadder_128 c_num_34(.data_in(dot_col_34), .sum(check_col_34));
bitsadder_128 c_num_35(.data_in(dot_col_35), .sum(check_col_35));
bitsadder_128 c_num_36(.data_in(dot_col_36), .sum(check_col_36));
bitsadder_128 c_num_37(.data_in(dot_col_37), .sum(check_col_37));
bitsadder_128 c_num_38(.data_in(dot_col_38), .sum(check_col_38));
bitsadder_128 c_num_39(.data_in(dot_col_39), .sum(check_col_39));
bitsadder_128 c_num_40(.data_in(dot_col_40), .sum(check_col_40));
bitsadder_128 c_num_41(.data_in(dot_col_41), .sum(check_col_41));
bitsadder_128 c_num_42(.data_in(dot_col_42), .sum(check_col_42));
bitsadder_128 c_num_43(.data_in(dot_col_43), .sum(check_col_43));
bitsadder_128 c_num_44(.data_in(dot_col_44), .sum(check_col_44));
bitsadder_128 c_num_45(.data_in(dot_col_45), .sum(check_col_45));
bitsadder_128 c_num_46(.data_in(dot_col_46), .sum(check_col_46));
bitsadder_128 c_num_47(.data_in(dot_col_47), .sum(check_col_47));
bitsadder_128 c_num_48(.data_in(dot_col_48), .sum(check_col_48));
bitsadder_128 c_num_49(.data_in(dot_col_49), .sum(check_col_49));
bitsadder_128 c_num_50(.data_in(dot_col_50), .sum(check_col_50));
bitsadder_128 c_num_51(.data_in(dot_col_51), .sum(check_col_51));
bitsadder_128 c_num_52(.data_in(dot_col_52), .sum(check_col_52));
bitsadder_128 c_num_53(.data_in(dot_col_53), .sum(check_col_53));
bitsadder_128 c_num_54(.data_in(dot_col_54), .sum(check_col_54));
bitsadder_128 c_num_55(.data_in(dot_col_55), .sum(check_col_55));
bitsadder_128 c_num_56(.data_in(dot_col_56), .sum(check_col_56));
bitsadder_128 c_num_57(.data_in(dot_col_57), .sum(check_col_57));
bitsadder_128 c_num_58(.data_in(dot_col_58), .sum(check_col_58));
bitsadder_128 c_num_59(.data_in(dot_col_59), .sum(check_col_59));
bitsadder_128 c_num_60(.data_in(dot_col_60), .sum(check_col_60));
bitsadder_128 c_num_61(.data_in(dot_col_61), .sum(check_col_61));
bitsadder_128 c_num_62(.data_in(dot_col_62), .sum(check_col_62));
bitsadder_128 c_num_63(.data_in(dot_col_63), .sum(check_col_63));
bitsadder_128 c_num_64(.data_in(dot_col_64), .sum(check_col_64));
bitsadder_128 c_num_65(.data_in(dot_col_65), .sum(check_col_65));
bitsadder_128 c_num_66(.data_in(dot_col_66), .sum(check_col_66));
bitsadder_128 c_num_67(.data_in(dot_col_67), .sum(check_col_67));
bitsadder_128 c_num_68(.data_in(dot_col_68), .sum(check_col_68));
bitsadder_128 c_num_69(.data_in(dot_col_69), .sum(check_col_69));
bitsadder_128 c_num_70(.data_in(dot_col_70), .sum(check_col_70));
bitsadder_128 c_num_71(.data_in(dot_col_71), .sum(check_col_71));
bitsadder_128 c_num_72(.data_in(dot_col_72), .sum(check_col_72));
bitsadder_128 c_num_73(.data_in(dot_col_73), .sum(check_col_73));
bitsadder_128 c_num_74(.data_in(dot_col_74), .sum(check_col_74));
bitsadder_128 c_num_75(.data_in(dot_col_75), .sum(check_col_75));
bitsadder_128 c_num_76(.data_in(dot_col_76), .sum(check_col_76));
bitsadder_128 c_num_77(.data_in(dot_col_77), .sum(check_col_77));
bitsadder_128 c_num_78(.data_in(dot_col_78), .sum(check_col_78));
bitsadder_128 c_num_79(.data_in(dot_col_79), .sum(check_col_79));
bitsadder_128 c_num_80(.data_in(dot_col_80), .sum(check_col_80));
bitsadder_128 c_num_81(.data_in(dot_col_81), .sum(check_col_81));
bitsadder_128 c_num_82(.data_in(dot_col_82), .sum(check_col_82));
bitsadder_128 c_num_83(.data_in(dot_col_83), .sum(check_col_83));
bitsadder_128 c_num_84(.data_in(dot_col_84), .sum(check_col_84));
bitsadder_128 c_num_85(.data_in(dot_col_85), .sum(check_col_85));
bitsadder_128 c_num_86(.data_in(dot_col_86), .sum(check_col_86));
bitsadder_128 c_num_87(.data_in(dot_col_87), .sum(check_col_87));
bitsadder_128 c_num_88(.data_in(dot_col_88), .sum(check_col_88));
bitsadder_128 c_num_89(.data_in(dot_col_89), .sum(check_col_89));
bitsadder_128 c_num_90(.data_in(dot_col_90), .sum(check_col_90));
bitsadder_128 c_num_91(.data_in(dot_col_91), .sum(check_col_91));
bitsadder_128 c_num_92(.data_in(dot_col_92), .sum(check_col_92));
bitsadder_128 c_num_93(.data_in(dot_col_93), .sum(check_col_93));
bitsadder_128 c_num_94(.data_in(dot_col_94), .sum(check_col_94));
bitsadder_128 c_num_95(.data_in(dot_col_95), .sum(check_col_95));
bitsadder_128 c_num_96(.data_in(dot_col_96), .sum(check_col_96));
bitsadder_128 c_num_97(.data_in(dot_col_97), .sum(check_col_97));
bitsadder_128 c_num_98(.data_in(dot_col_98), .sum(check_col_98));
bitsadder_128 c_num_99(.data_in(dot_col_99), .sum(check_col_99));
bitsadder_128 c_num_100(.data_in(dot_col_100), .sum(check_col_100));
bitsadder_128 c_num_101(.data_in(dot_col_101), .sum(check_col_101));
bitsadder_128 c_num_102(.data_in(dot_col_102), .sum(check_col_102));
bitsadder_128 c_num_103(.data_in(dot_col_103), .sum(check_col_103));
bitsadder_128 c_num_104(.data_in(dot_col_104), .sum(check_col_104));
bitsadder_128 c_num_105(.data_in(dot_col_105), .sum(check_col_105));
bitsadder_128 c_num_106(.data_in(dot_col_106), .sum(check_col_106));
bitsadder_128 c_num_107(.data_in(dot_col_107), .sum(check_col_107));
bitsadder_128 c_num_108(.data_in(dot_col_108), .sum(check_col_108));
bitsadder_128 c_num_109(.data_in(dot_col_109), .sum(check_col_109));
bitsadder_128 c_num_110(.data_in(dot_col_110), .sum(check_col_110));
bitsadder_128 c_num_111(.data_in(dot_col_111), .sum(check_col_111));
bitsadder_128 c_num_112(.data_in(dot_col_112), .sum(check_col_112));
bitsadder_128 c_num_113(.data_in(dot_col_113), .sum(check_col_113));
bitsadder_128 c_num_114(.data_in(dot_col_114), .sum(check_col_114));
bitsadder_128 c_num_115(.data_in(dot_col_115), .sum(check_col_115));
bitsadder_128 c_num_116(.data_in(dot_col_116), .sum(check_col_116));
bitsadder_128 c_num_117(.data_in(dot_col_117), .sum(check_col_117));
bitsadder_128 c_num_118(.data_in(dot_col_118), .sum(check_col_118));
bitsadder_128 c_num_119(.data_in(dot_col_119), .sum(check_col_119));
bitsadder_128 c_num_120(.data_in(dot_col_120), .sum(check_col_120));
bitsadder_128 c_num_121(.data_in(dot_col_121), .sum(check_col_121));
bitsadder_128 c_num_122(.data_in(dot_col_122), .sum(check_col_122));
bitsadder_128 c_num_123(.data_in(dot_col_123), .sum(check_col_123));
bitsadder_128 c_num_124(.data_in(dot_col_124), .sum(check_col_124));
bitsadder_128 c_num_125(.data_in(dot_col_125), .sum(check_col_125));
bitsadder_128 c_num_126(.data_in(dot_col_126), .sum(check_col_126));
bitsadder_128 c_num_127(.data_in(dot_col_127), .sum(check_col_127));
bitsadder_128 c_num_128(.data_in(dot_col_128), .sum(check_col_128));
bitsadder_128 c_num_129(.data_in(dot_col_129), .sum(check_col_129));
bitsadder_128 c_num_130(.data_in(dot_col_130), .sum(check_col_130));
bitsadder_128 c_num_131(.data_in(dot_col_131), .sum(check_col_131));
bitsadder_128 c_num_132(.data_in(dot_col_132), .sum(check_col_132));
bitsadder_128 c_num_133(.data_in(dot_col_133), .sum(check_col_133));
bitsadder_128 c_num_134(.data_in(dot_col_134), .sum(check_col_134));
bitsadder_128 c_num_135(.data_in(dot_col_135), .sum(check_col_135));
bitsadder_128 c_num_136(.data_in(dot_col_136), .sum(check_col_136));
bitsadder_128 c_num_137(.data_in(dot_col_137), .sum(check_col_137));
bitsadder_128 c_num_138(.data_in(dot_col_138), .sum(check_col_138));
bitsadder_128 c_num_139(.data_in(dot_col_139), .sum(check_col_139));
bitsadder_128 c_num_140(.data_in(dot_col_140), .sum(check_col_140));
bitsadder_128 c_num_141(.data_in(dot_col_141), .sum(check_col_141));
bitsadder_128 c_num_142(.data_in(dot_col_142), .sum(check_col_142));
bitsadder_128 c_num_143(.data_in(dot_col_143), .sum(check_col_143));
bitsadder_128 c_num_144(.data_in(dot_col_144), .sum(check_col_144));
bitsadder_128 c_num_145(.data_in(dot_col_145), .sum(check_col_145));
bitsadder_128 c_num_146(.data_in(dot_col_146), .sum(check_col_146));
bitsadder_128 c_num_147(.data_in(dot_col_147), .sum(check_col_147));
bitsadder_128 c_num_148(.data_in(dot_col_148), .sum(check_col_148));
bitsadder_128 c_num_149(.data_in(dot_col_149), .sum(check_col_149));
bitsadder_128 c_num_150(.data_in(dot_col_150), .sum(check_col_150));
bitsadder_128 c_num_151(.data_in(dot_col_151), .sum(check_col_151));
bitsadder_128 c_num_152(.data_in(dot_col_152), .sum(check_col_152));
bitsadder_128 c_num_153(.data_in(dot_col_153), .sum(check_col_153));
bitsadder_128 c_num_154(.data_in(dot_col_154), .sum(check_col_154));
bitsadder_128 c_num_155(.data_in(dot_col_155), .sum(check_col_155));
bitsadder_128 c_num_156(.data_in(dot_col_156), .sum(check_col_156));
bitsadder_128 c_num_157(.data_in(dot_col_157), .sum(check_col_157));
bitsadder_128 c_num_158(.data_in(dot_col_158), .sum(check_col_158));
bitsadder_128 c_num_159(.data_in(dot_col_159), .sum(check_col_159));
bitsadder_128 c_num_160(.data_in(dot_col_160), .sum(check_col_160));
bitsadder_128 c_num_161(.data_in(dot_col_161), .sum(check_col_161));
bitsadder_128 c_num_162(.data_in(dot_col_162), .sum(check_col_162));
bitsadder_128 c_num_163(.data_in(dot_col_163), .sum(check_col_163));
bitsadder_128 c_num_164(.data_in(dot_col_164), .sum(check_col_164));
bitsadder_128 c_num_165(.data_in(dot_col_165), .sum(check_col_165));
bitsadder_128 c_num_166(.data_in(dot_col_166), .sum(check_col_166));
bitsadder_128 c_num_167(.data_in(dot_col_167), .sum(check_col_167));
bitsadder_128 c_num_168(.data_in(dot_col_168), .sum(check_col_168));
bitsadder_128 c_num_169(.data_in(dot_col_169), .sum(check_col_169));
bitsadder_128 c_num_170(.data_in(dot_col_170), .sum(check_col_170));
bitsadder_128 c_num_171(.data_in(dot_col_171), .sum(check_col_171));
bitsadder_128 c_num_172(.data_in(dot_col_172), .sum(check_col_172));
bitsadder_128 c_num_173(.data_in(dot_col_173), .sum(check_col_173));
bitsadder_128 c_num_174(.data_in(dot_col_174), .sum(check_col_174));
bitsadder_128 c_num_175(.data_in(dot_col_175), .sum(check_col_175));
bitsadder_128 c_num_176(.data_in(dot_col_176), .sum(check_col_176));
bitsadder_128 c_num_177(.data_in(dot_col_177), .sum(check_col_177));
bitsadder_128 c_num_178(.data_in(dot_col_178), .sum(check_col_178));
bitsadder_128 c_num_179(.data_in(dot_col_179), .sum(check_col_179));
bitsadder_128 c_num_180(.data_in(dot_col_180), .sum(check_col_180));
bitsadder_128 c_num_181(.data_in(dot_col_181), .sum(check_col_181));
bitsadder_128 c_num_182(.data_in(dot_col_182), .sum(check_col_182));
bitsadder_128 c_num_183(.data_in(dot_col_183), .sum(check_col_183));
bitsadder_128 c_num_184(.data_in(dot_col_184), .sum(check_col_184));
bitsadder_128 c_num_185(.data_in(dot_col_185), .sum(check_col_185));
bitsadder_128 c_num_186(.data_in(dot_col_186), .sum(check_col_186));
bitsadder_128 c_num_187(.data_in(dot_col_187), .sum(check_col_187));
bitsadder_128 c_num_188(.data_in(dot_col_188), .sum(check_col_188));
bitsadder_128 c_num_189(.data_in(dot_col_189), .sum(check_col_189));
bitsadder_128 c_num_190(.data_in(dot_col_190), .sum(check_col_190));
bitsadder_128 c_num_191(.data_in(dot_col_191), .sum(check_col_191));
bitsadder_128 c_num_192(.data_in(dot_col_192), .sum(check_col_192));
bitsadder_128 c_num_193(.data_in(dot_col_193), .sum(check_col_193));
bitsadder_128 c_num_194(.data_in(dot_col_194), .sum(check_col_194));
bitsadder_128 c_num_195(.data_in(dot_col_195), .sum(check_col_195));
bitsadder_128 c_num_196(.data_in(dot_col_196), .sum(check_col_196));
bitsadder_128 c_num_197(.data_in(dot_col_197), .sum(check_col_197));
bitsadder_128 c_num_198(.data_in(dot_col_198), .sum(check_col_198));
bitsadder_128 c_num_199(.data_in(dot_col_199), .sum(check_col_199));
bitsadder_128 c_num_200(.data_in(dot_col_200), .sum(check_col_200));
bitsadder_128 c_num_201(.data_in(dot_col_201), .sum(check_col_201));
bitsadder_128 c_num_202(.data_in(dot_col_202), .sum(check_col_202));
bitsadder_128 c_num_203(.data_in(dot_col_203), .sum(check_col_203));
bitsadder_128 c_num_204(.data_in(dot_col_204), .sum(check_col_204));
bitsadder_128 c_num_205(.data_in(dot_col_205), .sum(check_col_205));
bitsadder_128 c_num_206(.data_in(dot_col_206), .sum(check_col_206));
bitsadder_128 c_num_207(.data_in(dot_col_207), .sum(check_col_207));
bitsadder_128 c_num_208(.data_in(dot_col_208), .sum(check_col_208));
bitsadder_128 c_num_209(.data_in(dot_col_209), .sum(check_col_209));
bitsadder_128 c_num_210(.data_in(dot_col_210), .sum(check_col_210));
bitsadder_128 c_num_211(.data_in(dot_col_211), .sum(check_col_211));
bitsadder_128 c_num_212(.data_in(dot_col_212), .sum(check_col_212));
bitsadder_128 c_num_213(.data_in(dot_col_213), .sum(check_col_213));
bitsadder_128 c_num_214(.data_in(dot_col_214), .sum(check_col_214));
bitsadder_128 c_num_215(.data_in(dot_col_215), .sum(check_col_215));
bitsadder_128 c_num_216(.data_in(dot_col_216), .sum(check_col_216));
bitsadder_128 c_num_217(.data_in(dot_col_217), .sum(check_col_217));
bitsadder_128 c_num_218(.data_in(dot_col_218), .sum(check_col_218));
bitsadder_128 c_num_219(.data_in(dot_col_219), .sum(check_col_219));
bitsadder_128 c_num_220(.data_in(dot_col_220), .sum(check_col_220));
bitsadder_128 c_num_221(.data_in(dot_col_221), .sum(check_col_221));
bitsadder_128 c_num_222(.data_in(dot_col_222), .sum(check_col_222));
bitsadder_128 c_num_223(.data_in(dot_col_223), .sum(check_col_223));
bitsadder_128 c_num_224(.data_in(dot_col_224), .sum(check_col_224));
bitsadder_128 c_num_225(.data_in(dot_col_225), .sum(check_col_225));
bitsadder_128 c_num_226(.data_in(dot_col_226), .sum(check_col_226));
bitsadder_128 c_num_227(.data_in(dot_col_227), .sum(check_col_227));
bitsadder_128 c_num_228(.data_in(dot_col_228), .sum(check_col_228));
bitsadder_128 c_num_229(.data_in(dot_col_229), .sum(check_col_229));
bitsadder_128 c_num_230(.data_in(dot_col_230), .sum(check_col_230));
bitsadder_128 c_num_231(.data_in(dot_col_231), .sum(check_col_231));
bitsadder_128 c_num_232(.data_in(dot_col_232), .sum(check_col_232));
bitsadder_128 c_num_233(.data_in(dot_col_233), .sum(check_col_233));
bitsadder_128 c_num_234(.data_in(dot_col_234), .sum(check_col_234));
bitsadder_128 c_num_235(.data_in(dot_col_235), .sum(check_col_235));
bitsadder_128 c_num_236(.data_in(dot_col_236), .sum(check_col_236));
bitsadder_128 c_num_237(.data_in(dot_col_237), .sum(check_col_237));
bitsadder_128 c_num_238(.data_in(dot_col_238), .sum(check_col_238));
bitsadder_128 c_num_239(.data_in(dot_col_239), .sum(check_col_239));
bitsadder_128 c_num_240(.data_in(dot_col_240), .sum(check_col_240));
bitsadder_128 c_num_241(.data_in(dot_col_241), .sum(check_col_241));
bitsadder_128 c_num_242(.data_in(dot_col_242), .sum(check_col_242));
bitsadder_128 c_num_243(.data_in(dot_col_243), .sum(check_col_243));
bitsadder_128 c_num_244(.data_in(dot_col_244), .sum(check_col_244));
bitsadder_128 c_num_245(.data_in(dot_col_245), .sum(check_col_245));
bitsadder_128 c_num_246(.data_in(dot_col_246), .sum(check_col_246));
bitsadder_128 c_num_247(.data_in(dot_col_247), .sum(check_col_247));
bitsadder_128 c_num_248(.data_in(dot_col_248), .sum(check_col_248));
bitsadder_128 c_num_249(.data_in(dot_col_249), .sum(check_col_249));
bitsadder_128 c_num_250(.data_in(dot_col_250), .sum(check_col_250));
bitsadder_128 c_num_251(.data_in(dot_col_251), .sum(check_col_251));
bitsadder_128 c_num_252(.data_in(dot_col_252), .sum(check_col_252));
bitsadder_128 c_num_253(.data_in(dot_col_253), .sum(check_col_253));
bitsadder_128 c_num_254(.data_in(dot_col_254), .sum(check_col_254));
bitsadder_128 c_num_255(.data_in(dot_col_255), .sum(check_col_255));


bitsadder_128 w_num_0(.data_in(dot_col_0 & form_array), .sum(wrong_col_0));
bitsadder_128 w_num_1(.data_in(dot_col_1 & form_array), .sum(wrong_col_1));
bitsadder_128 w_num_2(.data_in(dot_col_2 & form_array), .sum(wrong_col_2));
bitsadder_128 w_num_3(.data_in(dot_col_3 & form_array), .sum(wrong_col_3));
bitsadder_128 w_num_4(.data_in(dot_col_4 & form_array), .sum(wrong_col_4));
bitsadder_128 w_num_5(.data_in(dot_col_5 & form_array), .sum(wrong_col_5));
bitsadder_128 w_num_6(.data_in(dot_col_6 & form_array), .sum(wrong_col_6));
bitsadder_128 w_num_7(.data_in(dot_col_7 & form_array), .sum(wrong_col_7));
bitsadder_128 w_num_8(.data_in(dot_col_8 & form_array), .sum(wrong_col_8));
bitsadder_128 w_num_9(.data_in(dot_col_9 & form_array), .sum(wrong_col_9));
bitsadder_128 w_num_10(.data_in(dot_col_10 & form_array), .sum(wrong_col_10));
bitsadder_128 w_num_11(.data_in(dot_col_11 & form_array), .sum(wrong_col_11));
bitsadder_128 w_num_12(.data_in(dot_col_12 & form_array), .sum(wrong_col_12));
bitsadder_128 w_num_13(.data_in(dot_col_13 & form_array), .sum(wrong_col_13));
bitsadder_128 w_num_14(.data_in(dot_col_14 & form_array), .sum(wrong_col_14));
bitsadder_128 w_num_15(.data_in(dot_col_15 & form_array), .sum(wrong_col_15));
bitsadder_128 w_num_16(.data_in(dot_col_16 & form_array), .sum(wrong_col_16));
bitsadder_128 w_num_17(.data_in(dot_col_17 & form_array), .sum(wrong_col_17));
bitsadder_128 w_num_18(.data_in(dot_col_18 & form_array), .sum(wrong_col_18));
bitsadder_128 w_num_19(.data_in(dot_col_19 & form_array), .sum(wrong_col_19));
bitsadder_128 w_num_20(.data_in(dot_col_20 & form_array), .sum(wrong_col_20));
bitsadder_128 w_num_21(.data_in(dot_col_21 & form_array), .sum(wrong_col_21));
bitsadder_128 w_num_22(.data_in(dot_col_22 & form_array), .sum(wrong_col_22));
bitsadder_128 w_num_23(.data_in(dot_col_23 & form_array), .sum(wrong_col_23));
bitsadder_128 w_num_24(.data_in(dot_col_24 & form_array), .sum(wrong_col_24));
bitsadder_128 w_num_25(.data_in(dot_col_25 & form_array), .sum(wrong_col_25));
bitsadder_128 w_num_26(.data_in(dot_col_26 & form_array), .sum(wrong_col_26));
bitsadder_128 w_num_27(.data_in(dot_col_27 & form_array), .sum(wrong_col_27));
bitsadder_128 w_num_28(.data_in(dot_col_28 & form_array), .sum(wrong_col_28));
bitsadder_128 w_num_29(.data_in(dot_col_29 & form_array), .sum(wrong_col_29));
bitsadder_128 w_num_30(.data_in(dot_col_30 & form_array), .sum(wrong_col_30));
bitsadder_128 w_num_31(.data_in(dot_col_31 & form_array), .sum(wrong_col_31));
bitsadder_128 w_num_32(.data_in(dot_col_32 & form_array), .sum(wrong_col_32));
bitsadder_128 w_num_33(.data_in(dot_col_33 & form_array), .sum(wrong_col_33));
bitsadder_128 w_num_34(.data_in(dot_col_34 & form_array), .sum(wrong_col_34));
bitsadder_128 w_num_35(.data_in(dot_col_35 & form_array), .sum(wrong_col_35));
bitsadder_128 w_num_36(.data_in(dot_col_36 & form_array), .sum(wrong_col_36));
bitsadder_128 w_num_37(.data_in(dot_col_37 & form_array), .sum(wrong_col_37));
bitsadder_128 w_num_38(.data_in(dot_col_38 & form_array), .sum(wrong_col_38));
bitsadder_128 w_num_39(.data_in(dot_col_39 & form_array), .sum(wrong_col_39));
bitsadder_128 w_num_40(.data_in(dot_col_40 & form_array), .sum(wrong_col_40));
bitsadder_128 w_num_41(.data_in(dot_col_41 & form_array), .sum(wrong_col_41));
bitsadder_128 w_num_42(.data_in(dot_col_42 & form_array), .sum(wrong_col_42));
bitsadder_128 w_num_43(.data_in(dot_col_43 & form_array), .sum(wrong_col_43));
bitsadder_128 w_num_44(.data_in(dot_col_44 & form_array), .sum(wrong_col_44));
bitsadder_128 w_num_45(.data_in(dot_col_45 & form_array), .sum(wrong_col_45));
bitsadder_128 w_num_46(.data_in(dot_col_46 & form_array), .sum(wrong_col_46));
bitsadder_128 w_num_47(.data_in(dot_col_47 & form_array), .sum(wrong_col_47));
bitsadder_128 w_num_48(.data_in(dot_col_48 & form_array), .sum(wrong_col_48));
bitsadder_128 w_num_49(.data_in(dot_col_49 & form_array), .sum(wrong_col_49));
bitsadder_128 w_num_50(.data_in(dot_col_50 & form_array), .sum(wrong_col_50));
bitsadder_128 w_num_51(.data_in(dot_col_51 & form_array), .sum(wrong_col_51));
bitsadder_128 w_num_52(.data_in(dot_col_52 & form_array), .sum(wrong_col_52));
bitsadder_128 w_num_53(.data_in(dot_col_53 & form_array), .sum(wrong_col_53));
bitsadder_128 w_num_54(.data_in(dot_col_54 & form_array), .sum(wrong_col_54));
bitsadder_128 w_num_55(.data_in(dot_col_55 & form_array), .sum(wrong_col_55));
bitsadder_128 w_num_56(.data_in(dot_col_56 & form_array), .sum(wrong_col_56));
bitsadder_128 w_num_57(.data_in(dot_col_57 & form_array), .sum(wrong_col_57));
bitsadder_128 w_num_58(.data_in(dot_col_58 & form_array), .sum(wrong_col_58));
bitsadder_128 w_num_59(.data_in(dot_col_59 & form_array), .sum(wrong_col_59));
bitsadder_128 w_num_60(.data_in(dot_col_60 & form_array), .sum(wrong_col_60));
bitsadder_128 w_num_61(.data_in(dot_col_61 & form_array), .sum(wrong_col_61));
bitsadder_128 w_num_62(.data_in(dot_col_62 & form_array), .sum(wrong_col_62));
bitsadder_128 w_num_63(.data_in(dot_col_63 & form_array), .sum(wrong_col_63));
bitsadder_128 w_num_64(.data_in(dot_col_64 & form_array), .sum(wrong_col_64));
bitsadder_128 w_num_65(.data_in(dot_col_65 & form_array), .sum(wrong_col_65));
bitsadder_128 w_num_66(.data_in(dot_col_66 & form_array), .sum(wrong_col_66));
bitsadder_128 w_num_67(.data_in(dot_col_67 & form_array), .sum(wrong_col_67));
bitsadder_128 w_num_68(.data_in(dot_col_68 & form_array), .sum(wrong_col_68));
bitsadder_128 w_num_69(.data_in(dot_col_69 & form_array), .sum(wrong_col_69));
bitsadder_128 w_num_70(.data_in(dot_col_70 & form_array), .sum(wrong_col_70));
bitsadder_128 w_num_71(.data_in(dot_col_71 & form_array), .sum(wrong_col_71));
bitsadder_128 w_num_72(.data_in(dot_col_72 & form_array), .sum(wrong_col_72));
bitsadder_128 w_num_73(.data_in(dot_col_73 & form_array), .sum(wrong_col_73));
bitsadder_128 w_num_74(.data_in(dot_col_74 & form_array), .sum(wrong_col_74));
bitsadder_128 w_num_75(.data_in(dot_col_75 & form_array), .sum(wrong_col_75));
bitsadder_128 w_num_76(.data_in(dot_col_76 & form_array), .sum(wrong_col_76));
bitsadder_128 w_num_77(.data_in(dot_col_77 & form_array), .sum(wrong_col_77));
bitsadder_128 w_num_78(.data_in(dot_col_78 & form_array), .sum(wrong_col_78));
bitsadder_128 w_num_79(.data_in(dot_col_79 & form_array), .sum(wrong_col_79));
bitsadder_128 w_num_80(.data_in(dot_col_80 & form_array), .sum(wrong_col_80));
bitsadder_128 w_num_81(.data_in(dot_col_81 & form_array), .sum(wrong_col_81));
bitsadder_128 w_num_82(.data_in(dot_col_82 & form_array), .sum(wrong_col_82));
bitsadder_128 w_num_83(.data_in(dot_col_83 & form_array), .sum(wrong_col_83));
bitsadder_128 w_num_84(.data_in(dot_col_84 & form_array), .sum(wrong_col_84));
bitsadder_128 w_num_85(.data_in(dot_col_85 & form_array), .sum(wrong_col_85));
bitsadder_128 w_num_86(.data_in(dot_col_86 & form_array), .sum(wrong_col_86));
bitsadder_128 w_num_87(.data_in(dot_col_87 & form_array), .sum(wrong_col_87));
bitsadder_128 w_num_88(.data_in(dot_col_88 & form_array), .sum(wrong_col_88));
bitsadder_128 w_num_89(.data_in(dot_col_89 & form_array), .sum(wrong_col_89));
bitsadder_128 w_num_90(.data_in(dot_col_90 & form_array), .sum(wrong_col_90));
bitsadder_128 w_num_91(.data_in(dot_col_91 & form_array), .sum(wrong_col_91));
bitsadder_128 w_num_92(.data_in(dot_col_92 & form_array), .sum(wrong_col_92));
bitsadder_128 w_num_93(.data_in(dot_col_93 & form_array), .sum(wrong_col_93));
bitsadder_128 w_num_94(.data_in(dot_col_94 & form_array), .sum(wrong_col_94));
bitsadder_128 w_num_95(.data_in(dot_col_95 & form_array), .sum(wrong_col_95));
bitsadder_128 w_num_96(.data_in(dot_col_96 & form_array), .sum(wrong_col_96));
bitsadder_128 w_num_97(.data_in(dot_col_97 & form_array), .sum(wrong_col_97));
bitsadder_128 w_num_98(.data_in(dot_col_98 & form_array), .sum(wrong_col_98));
bitsadder_128 w_num_99(.data_in(dot_col_99 & form_array), .sum(wrong_col_99));
bitsadder_128 w_num_100(.data_in(dot_col_100 & form_array), .sum(wrong_col_100));
bitsadder_128 w_num_101(.data_in(dot_col_101 & form_array), .sum(wrong_col_101));
bitsadder_128 w_num_102(.data_in(dot_col_102 & form_array), .sum(wrong_col_102));
bitsadder_128 w_num_103(.data_in(dot_col_103 & form_array), .sum(wrong_col_103));
bitsadder_128 w_num_104(.data_in(dot_col_104 & form_array), .sum(wrong_col_104));
bitsadder_128 w_num_105(.data_in(dot_col_105 & form_array), .sum(wrong_col_105));
bitsadder_128 w_num_106(.data_in(dot_col_106 & form_array), .sum(wrong_col_106));
bitsadder_128 w_num_107(.data_in(dot_col_107 & form_array), .sum(wrong_col_107));
bitsadder_128 w_num_108(.data_in(dot_col_108 & form_array), .sum(wrong_col_108));
bitsadder_128 w_num_109(.data_in(dot_col_109 & form_array), .sum(wrong_col_109));
bitsadder_128 w_num_110(.data_in(dot_col_110 & form_array), .sum(wrong_col_110));
bitsadder_128 w_num_111(.data_in(dot_col_111 & form_array), .sum(wrong_col_111));
bitsadder_128 w_num_112(.data_in(dot_col_112 & form_array), .sum(wrong_col_112));
bitsadder_128 w_num_113(.data_in(dot_col_113 & form_array), .sum(wrong_col_113));
bitsadder_128 w_num_114(.data_in(dot_col_114 & form_array), .sum(wrong_col_114));
bitsadder_128 w_num_115(.data_in(dot_col_115 & form_array), .sum(wrong_col_115));
bitsadder_128 w_num_116(.data_in(dot_col_116 & form_array), .sum(wrong_col_116));
bitsadder_128 w_num_117(.data_in(dot_col_117 & form_array), .sum(wrong_col_117));
bitsadder_128 w_num_118(.data_in(dot_col_118 & form_array), .sum(wrong_col_118));
bitsadder_128 w_num_119(.data_in(dot_col_119 & form_array), .sum(wrong_col_119));
bitsadder_128 w_num_120(.data_in(dot_col_120 & form_array), .sum(wrong_col_120));
bitsadder_128 w_num_121(.data_in(dot_col_121 & form_array), .sum(wrong_col_121));
bitsadder_128 w_num_122(.data_in(dot_col_122 & form_array), .sum(wrong_col_122));
bitsadder_128 w_num_123(.data_in(dot_col_123 & form_array), .sum(wrong_col_123));
bitsadder_128 w_num_124(.data_in(dot_col_124 & form_array), .sum(wrong_col_124));
bitsadder_128 w_num_125(.data_in(dot_col_125 & form_array), .sum(wrong_col_125));
bitsadder_128 w_num_126(.data_in(dot_col_126 & form_array), .sum(wrong_col_126));
bitsadder_128 w_num_127(.data_in(dot_col_127 & form_array), .sum(wrong_col_127));
bitsadder_128 w_num_128(.data_in(dot_col_128 & form_array), .sum(wrong_col_128));
bitsadder_128 w_num_129(.data_in(dot_col_129 & form_array), .sum(wrong_col_129));
bitsadder_128 w_num_130(.data_in(dot_col_130 & form_array), .sum(wrong_col_130));
bitsadder_128 w_num_131(.data_in(dot_col_131 & form_array), .sum(wrong_col_131));
bitsadder_128 w_num_132(.data_in(dot_col_132 & form_array), .sum(wrong_col_132));
bitsadder_128 w_num_133(.data_in(dot_col_133 & form_array), .sum(wrong_col_133));
bitsadder_128 w_num_134(.data_in(dot_col_134 & form_array), .sum(wrong_col_134));
bitsadder_128 w_num_135(.data_in(dot_col_135 & form_array), .sum(wrong_col_135));
bitsadder_128 w_num_136(.data_in(dot_col_136 & form_array), .sum(wrong_col_136));
bitsadder_128 w_num_137(.data_in(dot_col_137 & form_array), .sum(wrong_col_137));
bitsadder_128 w_num_138(.data_in(dot_col_138 & form_array), .sum(wrong_col_138));
bitsadder_128 w_num_139(.data_in(dot_col_139 & form_array), .sum(wrong_col_139));
bitsadder_128 w_num_140(.data_in(dot_col_140 & form_array), .sum(wrong_col_140));
bitsadder_128 w_num_141(.data_in(dot_col_141 & form_array), .sum(wrong_col_141));
bitsadder_128 w_num_142(.data_in(dot_col_142 & form_array), .sum(wrong_col_142));
bitsadder_128 w_num_143(.data_in(dot_col_143 & form_array), .sum(wrong_col_143));
bitsadder_128 w_num_144(.data_in(dot_col_144 & form_array), .sum(wrong_col_144));
bitsadder_128 w_num_145(.data_in(dot_col_145 & form_array), .sum(wrong_col_145));
bitsadder_128 w_num_146(.data_in(dot_col_146 & form_array), .sum(wrong_col_146));
bitsadder_128 w_num_147(.data_in(dot_col_147 & form_array), .sum(wrong_col_147));
bitsadder_128 w_num_148(.data_in(dot_col_148 & form_array), .sum(wrong_col_148));
bitsadder_128 w_num_149(.data_in(dot_col_149 & form_array), .sum(wrong_col_149));
bitsadder_128 w_num_150(.data_in(dot_col_150 & form_array), .sum(wrong_col_150));
bitsadder_128 w_num_151(.data_in(dot_col_151 & form_array), .sum(wrong_col_151));
bitsadder_128 w_num_152(.data_in(dot_col_152 & form_array), .sum(wrong_col_152));
bitsadder_128 w_num_153(.data_in(dot_col_153 & form_array), .sum(wrong_col_153));
bitsadder_128 w_num_154(.data_in(dot_col_154 & form_array), .sum(wrong_col_154));
bitsadder_128 w_num_155(.data_in(dot_col_155 & form_array), .sum(wrong_col_155));
bitsadder_128 w_num_156(.data_in(dot_col_156 & form_array), .sum(wrong_col_156));
bitsadder_128 w_num_157(.data_in(dot_col_157 & form_array), .sum(wrong_col_157));
bitsadder_128 w_num_158(.data_in(dot_col_158 & form_array), .sum(wrong_col_158));
bitsadder_128 w_num_159(.data_in(dot_col_159 & form_array), .sum(wrong_col_159));
bitsadder_128 w_num_160(.data_in(dot_col_160 & form_array), .sum(wrong_col_160));
bitsadder_128 w_num_161(.data_in(dot_col_161 & form_array), .sum(wrong_col_161));
bitsadder_128 w_num_162(.data_in(dot_col_162 & form_array), .sum(wrong_col_162));
bitsadder_128 w_num_163(.data_in(dot_col_163 & form_array), .sum(wrong_col_163));
bitsadder_128 w_num_164(.data_in(dot_col_164 & form_array), .sum(wrong_col_164));
bitsadder_128 w_num_165(.data_in(dot_col_165 & form_array), .sum(wrong_col_165));
bitsadder_128 w_num_166(.data_in(dot_col_166 & form_array), .sum(wrong_col_166));
bitsadder_128 w_num_167(.data_in(dot_col_167 & form_array), .sum(wrong_col_167));
bitsadder_128 w_num_168(.data_in(dot_col_168 & form_array), .sum(wrong_col_168));
bitsadder_128 w_num_169(.data_in(dot_col_169 & form_array), .sum(wrong_col_169));
bitsadder_128 w_num_170(.data_in(dot_col_170 & form_array), .sum(wrong_col_170));
bitsadder_128 w_num_171(.data_in(dot_col_171 & form_array), .sum(wrong_col_171));
bitsadder_128 w_num_172(.data_in(dot_col_172 & form_array), .sum(wrong_col_172));
bitsadder_128 w_num_173(.data_in(dot_col_173 & form_array), .sum(wrong_col_173));
bitsadder_128 w_num_174(.data_in(dot_col_174 & form_array), .sum(wrong_col_174));
bitsadder_128 w_num_175(.data_in(dot_col_175 & form_array), .sum(wrong_col_175));
bitsadder_128 w_num_176(.data_in(dot_col_176 & form_array), .sum(wrong_col_176));
bitsadder_128 w_num_177(.data_in(dot_col_177 & form_array), .sum(wrong_col_177));
bitsadder_128 w_num_178(.data_in(dot_col_178 & form_array), .sum(wrong_col_178));
bitsadder_128 w_num_179(.data_in(dot_col_179 & form_array), .sum(wrong_col_179));
bitsadder_128 w_num_180(.data_in(dot_col_180 & form_array), .sum(wrong_col_180));
bitsadder_128 w_num_181(.data_in(dot_col_181 & form_array), .sum(wrong_col_181));
bitsadder_128 w_num_182(.data_in(dot_col_182 & form_array), .sum(wrong_col_182));
bitsadder_128 w_num_183(.data_in(dot_col_183 & form_array), .sum(wrong_col_183));
bitsadder_128 w_num_184(.data_in(dot_col_184 & form_array), .sum(wrong_col_184));
bitsadder_128 w_num_185(.data_in(dot_col_185 & form_array), .sum(wrong_col_185));
bitsadder_128 w_num_186(.data_in(dot_col_186 & form_array), .sum(wrong_col_186));
bitsadder_128 w_num_187(.data_in(dot_col_187 & form_array), .sum(wrong_col_187));
bitsadder_128 w_num_188(.data_in(dot_col_188 & form_array), .sum(wrong_col_188));
bitsadder_128 w_num_189(.data_in(dot_col_189 & form_array), .sum(wrong_col_189));
bitsadder_128 w_num_190(.data_in(dot_col_190 & form_array), .sum(wrong_col_190));
bitsadder_128 w_num_191(.data_in(dot_col_191 & form_array), .sum(wrong_col_191));
bitsadder_128 w_num_192(.data_in(dot_col_192 & form_array), .sum(wrong_col_192));
bitsadder_128 w_num_193(.data_in(dot_col_193 & form_array), .sum(wrong_col_193));
bitsadder_128 w_num_194(.data_in(dot_col_194 & form_array), .sum(wrong_col_194));
bitsadder_128 w_num_195(.data_in(dot_col_195 & form_array), .sum(wrong_col_195));
bitsadder_128 w_num_196(.data_in(dot_col_196 & form_array), .sum(wrong_col_196));
bitsadder_128 w_num_197(.data_in(dot_col_197 & form_array), .sum(wrong_col_197));
bitsadder_128 w_num_198(.data_in(dot_col_198 & form_array), .sum(wrong_col_198));
bitsadder_128 w_num_199(.data_in(dot_col_199 & form_array), .sum(wrong_col_199));
bitsadder_128 w_num_200(.data_in(dot_col_200 & form_array), .sum(wrong_col_200));
bitsadder_128 w_num_201(.data_in(dot_col_201 & form_array), .sum(wrong_col_201));
bitsadder_128 w_num_202(.data_in(dot_col_202 & form_array), .sum(wrong_col_202));
bitsadder_128 w_num_203(.data_in(dot_col_203 & form_array), .sum(wrong_col_203));
bitsadder_128 w_num_204(.data_in(dot_col_204 & form_array), .sum(wrong_col_204));
bitsadder_128 w_num_205(.data_in(dot_col_205 & form_array), .sum(wrong_col_205));
bitsadder_128 w_num_206(.data_in(dot_col_206 & form_array), .sum(wrong_col_206));
bitsadder_128 w_num_207(.data_in(dot_col_207 & form_array), .sum(wrong_col_207));
bitsadder_128 w_num_208(.data_in(dot_col_208 & form_array), .sum(wrong_col_208));
bitsadder_128 w_num_209(.data_in(dot_col_209 & form_array), .sum(wrong_col_209));
bitsadder_128 w_num_210(.data_in(dot_col_210 & form_array), .sum(wrong_col_210));
bitsadder_128 w_num_211(.data_in(dot_col_211 & form_array), .sum(wrong_col_211));
bitsadder_128 w_num_212(.data_in(dot_col_212 & form_array), .sum(wrong_col_212));
bitsadder_128 w_num_213(.data_in(dot_col_213 & form_array), .sum(wrong_col_213));
bitsadder_128 w_num_214(.data_in(dot_col_214 & form_array), .sum(wrong_col_214));
bitsadder_128 w_num_215(.data_in(dot_col_215 & form_array), .sum(wrong_col_215));
bitsadder_128 w_num_216(.data_in(dot_col_216 & form_array), .sum(wrong_col_216));
bitsadder_128 w_num_217(.data_in(dot_col_217 & form_array), .sum(wrong_col_217));
bitsadder_128 w_num_218(.data_in(dot_col_218 & form_array), .sum(wrong_col_218));
bitsadder_128 w_num_219(.data_in(dot_col_219 & form_array), .sum(wrong_col_219));
bitsadder_128 w_num_220(.data_in(dot_col_220 & form_array), .sum(wrong_col_220));
bitsadder_128 w_num_221(.data_in(dot_col_221 & form_array), .sum(wrong_col_221));
bitsadder_128 w_num_222(.data_in(dot_col_222 & form_array), .sum(wrong_col_222));
bitsadder_128 w_num_223(.data_in(dot_col_223 & form_array), .sum(wrong_col_223));
bitsadder_128 w_num_224(.data_in(dot_col_224 & form_array), .sum(wrong_col_224));
bitsadder_128 w_num_225(.data_in(dot_col_225 & form_array), .sum(wrong_col_225));
bitsadder_128 w_num_226(.data_in(dot_col_226 & form_array), .sum(wrong_col_226));
bitsadder_128 w_num_227(.data_in(dot_col_227 & form_array), .sum(wrong_col_227));
bitsadder_128 w_num_228(.data_in(dot_col_228 & form_array), .sum(wrong_col_228));
bitsadder_128 w_num_229(.data_in(dot_col_229 & form_array), .sum(wrong_col_229));
bitsadder_128 w_num_230(.data_in(dot_col_230 & form_array), .sum(wrong_col_230));
bitsadder_128 w_num_231(.data_in(dot_col_231 & form_array), .sum(wrong_col_231));
bitsadder_128 w_num_232(.data_in(dot_col_232 & form_array), .sum(wrong_col_232));
bitsadder_128 w_num_233(.data_in(dot_col_233 & form_array), .sum(wrong_col_233));
bitsadder_128 w_num_234(.data_in(dot_col_234 & form_array), .sum(wrong_col_234));
bitsadder_128 w_num_235(.data_in(dot_col_235 & form_array), .sum(wrong_col_235));
bitsadder_128 w_num_236(.data_in(dot_col_236 & form_array), .sum(wrong_col_236));
bitsadder_128 w_num_237(.data_in(dot_col_237 & form_array), .sum(wrong_col_237));
bitsadder_128 w_num_238(.data_in(dot_col_238 & form_array), .sum(wrong_col_238));
bitsadder_128 w_num_239(.data_in(dot_col_239 & form_array), .sum(wrong_col_239));
bitsadder_128 w_num_240(.data_in(dot_col_240 & form_array), .sum(wrong_col_240));
bitsadder_128 w_num_241(.data_in(dot_col_241 & form_array), .sum(wrong_col_241));
bitsadder_128 w_num_242(.data_in(dot_col_242 & form_array), .sum(wrong_col_242));
bitsadder_128 w_num_243(.data_in(dot_col_243 & form_array), .sum(wrong_col_243));
bitsadder_128 w_num_244(.data_in(dot_col_244 & form_array), .sum(wrong_col_244));
bitsadder_128 w_num_245(.data_in(dot_col_245 & form_array), .sum(wrong_col_245));
bitsadder_128 w_num_246(.data_in(dot_col_246 & form_array), .sum(wrong_col_246));
bitsadder_128 w_num_247(.data_in(dot_col_247 & form_array), .sum(wrong_col_247));
bitsadder_128 w_num_248(.data_in(dot_col_248 & form_array), .sum(wrong_col_248));
bitsadder_128 w_num_249(.data_in(dot_col_249 & form_array), .sum(wrong_col_249));
bitsadder_128 w_num_250(.data_in(dot_col_250 & form_array), .sum(wrong_col_250));
bitsadder_128 w_num_251(.data_in(dot_col_251 & form_array), .sum(wrong_col_251));
bitsadder_128 w_num_252(.data_in(dot_col_252 & form_array), .sum(wrong_col_252));
bitsadder_128 w_num_253(.data_in(dot_col_253 & form_array), .sum(wrong_col_253));
bitsadder_128 w_num_254(.data_in(dot_col_254 & form_array), .sum(wrong_col_254));
bitsadder_128 w_num_255(.data_in(dot_col_255 & form_array), .sum(wrong_col_255));


//Edit code:

always@(posedge clk or negedge rst) begin
if(!rst) begin
state <= init;
free_flag <= 1'b0;
valid_flag <= 1'b0;
iter_flag <= 1'b0;
iter_cnt <= 'd0;
deout_reg <= 'd0;
end
else begin

case(state)

init: begin
free_flag <= 1'b1;
tx_buffer <= 'd0;
form_array <= 'd0;
state <= getin;

end


getin: begin
if(work) begin
    tx_buffer <= tx;
    update_buffer <= tx;
    free_flag <= 1'b0;
    valid_flag <= 1'b0;
    iter_flag <= 1'b1;
    deout_reg <= 'd0;
    state <= dot;
end
else begin
    if (iter_flag) begin
        tx_buffer <= update_buffer;
        state <= dot;
    end
    else begin
        state <= getin;
    end
end

end


dot: begin
integer i;
for(i=0;i<256;i=i+1) begin
    dotarray[i] <= Harray[i] & tx_buffer;
end
state <= judge;

end


judge: begin
form_array <= row_sum_lastbit;
if(form_array == 'd0) begin
    state <= decode;
end
else begin
    valid_flag <= 1'b0;
    state <= check;
end

end


check: begin

check_cnt[0] <= ((check_col_0) >> 1);
check_cnt[1] <= ((check_col_1) >> 1);
check_cnt[2] <= ((check_col_2) >> 1);
check_cnt[3] <= ((check_col_3) >> 1);
check_cnt[4] <= ((check_col_4) >> 1);
check_cnt[5] <= ((check_col_5) >> 1);
check_cnt[6] <= ((check_col_6) >> 1);
check_cnt[7] <= ((check_col_7) >> 1);
check_cnt[8] <= ((check_col_8) >> 1);
check_cnt[9] <= ((check_col_9) >> 1);
check_cnt[10] <= ((check_col_10) >> 1);
check_cnt[11] <= ((check_col_11) >> 1);
check_cnt[12] <= ((check_col_12) >> 1);
check_cnt[13] <= ((check_col_13) >> 1);
check_cnt[14] <= ((check_col_14) >> 1);
check_cnt[15] <= ((check_col_15) >> 1);
check_cnt[16] <= ((check_col_16) >> 1);
check_cnt[17] <= ((check_col_17) >> 1);
check_cnt[18] <= ((check_col_18) >> 1);
check_cnt[19] <= ((check_col_19) >> 1);
check_cnt[20] <= ((check_col_20) >> 1);
check_cnt[21] <= ((check_col_21) >> 1);
check_cnt[22] <= ((check_col_22) >> 1);
check_cnt[23] <= ((check_col_23) >> 1);
check_cnt[24] <= ((check_col_24) >> 1);
check_cnt[25] <= ((check_col_25) >> 1);
check_cnt[26] <= ((check_col_26) >> 1);
check_cnt[27] <= ((check_col_27) >> 1);
check_cnt[28] <= ((check_col_28) >> 1);
check_cnt[29] <= ((check_col_29) >> 1);
check_cnt[30] <= ((check_col_30) >> 1);
check_cnt[31] <= ((check_col_31) >> 1);
check_cnt[32] <= ((check_col_32) >> 1);
check_cnt[33] <= ((check_col_33) >> 1);
check_cnt[34] <= ((check_col_34) >> 1);
check_cnt[35] <= ((check_col_35) >> 1);
check_cnt[36] <= ((check_col_36) >> 1);
check_cnt[37] <= ((check_col_37) >> 1);
check_cnt[38] <= ((check_col_38) >> 1);
check_cnt[39] <= ((check_col_39) >> 1);
check_cnt[40] <= ((check_col_40) >> 1);
check_cnt[41] <= ((check_col_41) >> 1);
check_cnt[42] <= ((check_col_42) >> 1);
check_cnt[43] <= ((check_col_43) >> 1);
check_cnt[44] <= ((check_col_44) >> 1);
check_cnt[45] <= ((check_col_45) >> 1);
check_cnt[46] <= ((check_col_46) >> 1);
check_cnt[47] <= ((check_col_47) >> 1);
check_cnt[48] <= ((check_col_48) >> 1);
check_cnt[49] <= ((check_col_49) >> 1);
check_cnt[50] <= ((check_col_50) >> 1);
check_cnt[51] <= ((check_col_51) >> 1);
check_cnt[52] <= ((check_col_52) >> 1);
check_cnt[53] <= ((check_col_53) >> 1);
check_cnt[54] <= ((check_col_54) >> 1);
check_cnt[55] <= ((check_col_55) >> 1);
check_cnt[56] <= ((check_col_56) >> 1);
check_cnt[57] <= ((check_col_57) >> 1);
check_cnt[58] <= ((check_col_58) >> 1);
check_cnt[59] <= ((check_col_59) >> 1);
check_cnt[60] <= ((check_col_60) >> 1);
check_cnt[61] <= ((check_col_61) >> 1);
check_cnt[62] <= ((check_col_62) >> 1);
check_cnt[63] <= ((check_col_63) >> 1);
check_cnt[64] <= ((check_col_64) >> 1);
check_cnt[65] <= ((check_col_65) >> 1);
check_cnt[66] <= ((check_col_66) >> 1);
check_cnt[67] <= ((check_col_67) >> 1);
check_cnt[68] <= ((check_col_68) >> 1);
check_cnt[69] <= ((check_col_69) >> 1);
check_cnt[70] <= ((check_col_70) >> 1);
check_cnt[71] <= ((check_col_71) >> 1);
check_cnt[72] <= ((check_col_72) >> 1);
check_cnt[73] <= ((check_col_73) >> 1);
check_cnt[74] <= ((check_col_74) >> 1);
check_cnt[75] <= ((check_col_75) >> 1);
check_cnt[76] <= ((check_col_76) >> 1);
check_cnt[77] <= ((check_col_77) >> 1);
check_cnt[78] <= ((check_col_78) >> 1);
check_cnt[79] <= ((check_col_79) >> 1);
check_cnt[80] <= ((check_col_80) >> 1);
check_cnt[81] <= ((check_col_81) >> 1);
check_cnt[82] <= ((check_col_82) >> 1);
check_cnt[83] <= ((check_col_83) >> 1);
check_cnt[84] <= ((check_col_84) >> 1);
check_cnt[85] <= ((check_col_85) >> 1);
check_cnt[86] <= ((check_col_86) >> 1);
check_cnt[87] <= ((check_col_87) >> 1);
check_cnt[88] <= ((check_col_88) >> 1);
check_cnt[89] <= ((check_col_89) >> 1);
check_cnt[90] <= ((check_col_90) >> 1);
check_cnt[91] <= ((check_col_91) >> 1);
check_cnt[92] <= ((check_col_92) >> 1);
check_cnt[93] <= ((check_col_93) >> 1);
check_cnt[94] <= ((check_col_94) >> 1);
check_cnt[95] <= ((check_col_95) >> 1);
check_cnt[96] <= ((check_col_96) >> 1);
check_cnt[97] <= ((check_col_97) >> 1);
check_cnt[98] <= ((check_col_98) >> 1);
check_cnt[99] <= ((check_col_99) >> 1);
check_cnt[100] <= ((check_col_100) >> 1);
check_cnt[101] <= ((check_col_101) >> 1);
check_cnt[102] <= ((check_col_102) >> 1);
check_cnt[103] <= ((check_col_103) >> 1);
check_cnt[104] <= ((check_col_104) >> 1);
check_cnt[105] <= ((check_col_105) >> 1);
check_cnt[106] <= ((check_col_106) >> 1);
check_cnt[107] <= ((check_col_107) >> 1);
check_cnt[108] <= ((check_col_108) >> 1);
check_cnt[109] <= ((check_col_109) >> 1);
check_cnt[110] <= ((check_col_110) >> 1);
check_cnt[111] <= ((check_col_111) >> 1);
check_cnt[112] <= ((check_col_112) >> 1);
check_cnt[113] <= ((check_col_113) >> 1);
check_cnt[114] <= ((check_col_114) >> 1);
check_cnt[115] <= ((check_col_115) >> 1);
check_cnt[116] <= ((check_col_116) >> 1);
check_cnt[117] <= ((check_col_117) >> 1);
check_cnt[118] <= ((check_col_118) >> 1);
check_cnt[119] <= ((check_col_119) >> 1);
check_cnt[120] <= ((check_col_120) >> 1);
check_cnt[121] <= ((check_col_121) >> 1);
check_cnt[122] <= ((check_col_122) >> 1);
check_cnt[123] <= ((check_col_123) >> 1);
check_cnt[124] <= ((check_col_124) >> 1);
check_cnt[125] <= ((check_col_125) >> 1);
check_cnt[126] <= ((check_col_126) >> 1);
check_cnt[127] <= ((check_col_127) >> 1);
check_cnt[128] <= ((check_col_128) >> 1);
check_cnt[129] <= ((check_col_129) >> 1);
check_cnt[130] <= ((check_col_130) >> 1);
check_cnt[131] <= ((check_col_131) >> 1);
check_cnt[132] <= ((check_col_132) >> 1);
check_cnt[133] <= ((check_col_133) >> 1);
check_cnt[134] <= ((check_col_134) >> 1);
check_cnt[135] <= ((check_col_135) >> 1);
check_cnt[136] <= ((check_col_136) >> 1);
check_cnt[137] <= ((check_col_137) >> 1);
check_cnt[138] <= ((check_col_138) >> 1);
check_cnt[139] <= ((check_col_139) >> 1);
check_cnt[140] <= ((check_col_140) >> 1);
check_cnt[141] <= ((check_col_141) >> 1);
check_cnt[142] <= ((check_col_142) >> 1);
check_cnt[143] <= ((check_col_143) >> 1);
check_cnt[144] <= ((check_col_144) >> 1);
check_cnt[145] <= ((check_col_145) >> 1);
check_cnt[146] <= ((check_col_146) >> 1);
check_cnt[147] <= ((check_col_147) >> 1);
check_cnt[148] <= ((check_col_148) >> 1);
check_cnt[149] <= ((check_col_149) >> 1);
check_cnt[150] <= ((check_col_150) >> 1);
check_cnt[151] <= ((check_col_151) >> 1);
check_cnt[152] <= ((check_col_152) >> 1);
check_cnt[153] <= ((check_col_153) >> 1);
check_cnt[154] <= ((check_col_154) >> 1);
check_cnt[155] <= ((check_col_155) >> 1);
check_cnt[156] <= ((check_col_156) >> 1);
check_cnt[157] <= ((check_col_157) >> 1);
check_cnt[158] <= ((check_col_158) >> 1);
check_cnt[159] <= ((check_col_159) >> 1);
check_cnt[160] <= ((check_col_160) >> 1);
check_cnt[161] <= ((check_col_161) >> 1);
check_cnt[162] <= ((check_col_162) >> 1);
check_cnt[163] <= ((check_col_163) >> 1);
check_cnt[164] <= ((check_col_164) >> 1);
check_cnt[165] <= ((check_col_165) >> 1);
check_cnt[166] <= ((check_col_166) >> 1);
check_cnt[167] <= ((check_col_167) >> 1);
check_cnt[168] <= ((check_col_168) >> 1);
check_cnt[169] <= ((check_col_169) >> 1);
check_cnt[170] <= ((check_col_170) >> 1);
check_cnt[171] <= ((check_col_171) >> 1);
check_cnt[172] <= ((check_col_172) >> 1);
check_cnt[173] <= ((check_col_173) >> 1);
check_cnt[174] <= ((check_col_174) >> 1);
check_cnt[175] <= ((check_col_175) >> 1);
check_cnt[176] <= ((check_col_176) >> 1);
check_cnt[177] <= ((check_col_177) >> 1);
check_cnt[178] <= ((check_col_178) >> 1);
check_cnt[179] <= ((check_col_179) >> 1);
check_cnt[180] <= ((check_col_180) >> 1);
check_cnt[181] <= ((check_col_181) >> 1);
check_cnt[182] <= ((check_col_182) >> 1);
check_cnt[183] <= ((check_col_183) >> 1);
check_cnt[184] <= ((check_col_184) >> 1);
check_cnt[185] <= ((check_col_185) >> 1);
check_cnt[186] <= ((check_col_186) >> 1);
check_cnt[187] <= ((check_col_187) >> 1);
check_cnt[188] <= ((check_col_188) >> 1);
check_cnt[189] <= ((check_col_189) >> 1);
check_cnt[190] <= ((check_col_190) >> 1);
check_cnt[191] <= ((check_col_191) >> 1);
check_cnt[192] <= ((check_col_192) >> 1);
check_cnt[193] <= ((check_col_193) >> 1);
check_cnt[194] <= ((check_col_194) >> 1);
check_cnt[195] <= ((check_col_195) >> 1);
check_cnt[196] <= ((check_col_196) >> 1);
check_cnt[197] <= ((check_col_197) >> 1);
check_cnt[198] <= ((check_col_198) >> 1);
check_cnt[199] <= ((check_col_199) >> 1);
check_cnt[200] <= ((check_col_200) >> 1);
check_cnt[201] <= ((check_col_201) >> 1);
check_cnt[202] <= ((check_col_202) >> 1);
check_cnt[203] <= ((check_col_203) >> 1);
check_cnt[204] <= ((check_col_204) >> 1);
check_cnt[205] <= ((check_col_205) >> 1);
check_cnt[206] <= ((check_col_206) >> 1);
check_cnt[207] <= ((check_col_207) >> 1);
check_cnt[208] <= ((check_col_208) >> 1);
check_cnt[209] <= ((check_col_209) >> 1);
check_cnt[210] <= ((check_col_210) >> 1);
check_cnt[211] <= ((check_col_211) >> 1);
check_cnt[212] <= ((check_col_212) >> 1);
check_cnt[213] <= ((check_col_213) >> 1);
check_cnt[214] <= ((check_col_214) >> 1);
check_cnt[215] <= ((check_col_215) >> 1);
check_cnt[216] <= ((check_col_216) >> 1);
check_cnt[217] <= ((check_col_217) >> 1);
check_cnt[218] <= ((check_col_218) >> 1);
check_cnt[219] <= ((check_col_219) >> 1);
check_cnt[220] <= ((check_col_220) >> 1);
check_cnt[221] <= ((check_col_221) >> 1);
check_cnt[222] <= ((check_col_222) >> 1);
check_cnt[223] <= ((check_col_223) >> 1);
check_cnt[224] <= ((check_col_224) >> 1);
check_cnt[225] <= ((check_col_225) >> 1);
check_cnt[226] <= ((check_col_226) >> 1);
check_cnt[227] <= ((check_col_227) >> 1);
check_cnt[228] <= ((check_col_228) >> 1);
check_cnt[229] <= ((check_col_229) >> 1);
check_cnt[230] <= ((check_col_230) >> 1);
check_cnt[231] <= ((check_col_231) >> 1);
check_cnt[232] <= ((check_col_232) >> 1);
check_cnt[233] <= ((check_col_233) >> 1);
check_cnt[234] <= ((check_col_234) >> 1);
check_cnt[235] <= ((check_col_235) >> 1);
check_cnt[236] <= ((check_col_236) >> 1);
check_cnt[237] <= ((check_col_237) >> 1);
check_cnt[238] <= ((check_col_238) >> 1);
check_cnt[239] <= ((check_col_239) >> 1);
check_cnt[240] <= ((check_col_240) >> 1);
check_cnt[241] <= ((check_col_241) >> 1);
check_cnt[242] <= ((check_col_242) >> 1);
check_cnt[243] <= ((check_col_243) >> 1);
check_cnt[244] <= ((check_col_244) >> 1);
check_cnt[245] <= ((check_col_245) >> 1);
check_cnt[246] <= ((check_col_246) >> 1);
check_cnt[247] <= ((check_col_247) >> 1);
check_cnt[248] <= ((check_col_248) >> 1);
check_cnt[249] <= ((check_col_249) >> 1);
check_cnt[250] <= ((check_col_250) >> 1);
check_cnt[251] <= ((check_col_251) >> 1);
check_cnt[252] <= ((check_col_252) >> 1);
check_cnt[253] <= ((check_col_253) >> 1);
check_cnt[254] <= ((check_col_254) >> 1);
check_cnt[255] <= ((check_col_255) >> 1);

wrong_cnt[0] <= wrong_col_0;
wrong_cnt[1] <= wrong_col_1;
wrong_cnt[2] <= wrong_col_2;
wrong_cnt[3] <= wrong_col_3;
wrong_cnt[4] <= wrong_col_4;
wrong_cnt[5] <= wrong_col_5;
wrong_cnt[6] <= wrong_col_6;
wrong_cnt[7] <= wrong_col_7;
wrong_cnt[8] <= wrong_col_8;
wrong_cnt[9] <= wrong_col_9;
wrong_cnt[10] <= wrong_col_10;
wrong_cnt[11] <= wrong_col_11;
wrong_cnt[12] <= wrong_col_12;
wrong_cnt[13] <= wrong_col_13;
wrong_cnt[14] <= wrong_col_14;
wrong_cnt[15] <= wrong_col_15;
wrong_cnt[16] <= wrong_col_16;
wrong_cnt[17] <= wrong_col_17;
wrong_cnt[18] <= wrong_col_18;
wrong_cnt[19] <= wrong_col_19;
wrong_cnt[20] <= wrong_col_20;
wrong_cnt[21] <= wrong_col_21;
wrong_cnt[22] <= wrong_col_22;
wrong_cnt[23] <= wrong_col_23;
wrong_cnt[24] <= wrong_col_24;
wrong_cnt[25] <= wrong_col_25;
wrong_cnt[26] <= wrong_col_26;
wrong_cnt[27] <= wrong_col_27;
wrong_cnt[28] <= wrong_col_28;
wrong_cnt[29] <= wrong_col_29;
wrong_cnt[30] <= wrong_col_30;
wrong_cnt[31] <= wrong_col_31;
wrong_cnt[32] <= wrong_col_32;
wrong_cnt[33] <= wrong_col_33;
wrong_cnt[34] <= wrong_col_34;
wrong_cnt[35] <= wrong_col_35;
wrong_cnt[36] <= wrong_col_36;
wrong_cnt[37] <= wrong_col_37;
wrong_cnt[38] <= wrong_col_38;
wrong_cnt[39] <= wrong_col_39;
wrong_cnt[40] <= wrong_col_40;
wrong_cnt[41] <= wrong_col_41;
wrong_cnt[42] <= wrong_col_42;
wrong_cnt[43] <= wrong_col_43;
wrong_cnt[44] <= wrong_col_44;
wrong_cnt[45] <= wrong_col_45;
wrong_cnt[46] <= wrong_col_46;
wrong_cnt[47] <= wrong_col_47;
wrong_cnt[48] <= wrong_col_48;
wrong_cnt[49] <= wrong_col_49;
wrong_cnt[50] <= wrong_col_50;
wrong_cnt[51] <= wrong_col_51;
wrong_cnt[52] <= wrong_col_52;
wrong_cnt[53] <= wrong_col_53;
wrong_cnt[54] <= wrong_col_54;
wrong_cnt[55] <= wrong_col_55;
wrong_cnt[56] <= wrong_col_56;
wrong_cnt[57] <= wrong_col_57;
wrong_cnt[58] <= wrong_col_58;
wrong_cnt[59] <= wrong_col_59;
wrong_cnt[60] <= wrong_col_60;
wrong_cnt[61] <= wrong_col_61;
wrong_cnt[62] <= wrong_col_62;
wrong_cnt[63] <= wrong_col_63;
wrong_cnt[64] <= wrong_col_64;
wrong_cnt[65] <= wrong_col_65;
wrong_cnt[66] <= wrong_col_66;
wrong_cnt[67] <= wrong_col_67;
wrong_cnt[68] <= wrong_col_68;
wrong_cnt[69] <= wrong_col_69;
wrong_cnt[70] <= wrong_col_70;
wrong_cnt[71] <= wrong_col_71;
wrong_cnt[72] <= wrong_col_72;
wrong_cnt[73] <= wrong_col_73;
wrong_cnt[74] <= wrong_col_74;
wrong_cnt[75] <= wrong_col_75;
wrong_cnt[76] <= wrong_col_76;
wrong_cnt[77] <= wrong_col_77;
wrong_cnt[78] <= wrong_col_78;
wrong_cnt[79] <= wrong_col_79;
wrong_cnt[80] <= wrong_col_80;
wrong_cnt[81] <= wrong_col_81;
wrong_cnt[82] <= wrong_col_82;
wrong_cnt[83] <= wrong_col_83;
wrong_cnt[84] <= wrong_col_84;
wrong_cnt[85] <= wrong_col_85;
wrong_cnt[86] <= wrong_col_86;
wrong_cnt[87] <= wrong_col_87;
wrong_cnt[88] <= wrong_col_88;
wrong_cnt[89] <= wrong_col_89;
wrong_cnt[90] <= wrong_col_90;
wrong_cnt[91] <= wrong_col_91;
wrong_cnt[92] <= wrong_col_92;
wrong_cnt[93] <= wrong_col_93;
wrong_cnt[94] <= wrong_col_94;
wrong_cnt[95] <= wrong_col_95;
wrong_cnt[96] <= wrong_col_96;
wrong_cnt[97] <= wrong_col_97;
wrong_cnt[98] <= wrong_col_98;
wrong_cnt[99] <= wrong_col_99;
wrong_cnt[100] <= wrong_col_100;
wrong_cnt[101] <= wrong_col_101;
wrong_cnt[102] <= wrong_col_102;
wrong_cnt[103] <= wrong_col_103;
wrong_cnt[104] <= wrong_col_104;
wrong_cnt[105] <= wrong_col_105;
wrong_cnt[106] <= wrong_col_106;
wrong_cnt[107] <= wrong_col_107;
wrong_cnt[108] <= wrong_col_108;
wrong_cnt[109] <= wrong_col_109;
wrong_cnt[110] <= wrong_col_110;
wrong_cnt[111] <= wrong_col_111;
wrong_cnt[112] <= wrong_col_112;
wrong_cnt[113] <= wrong_col_113;
wrong_cnt[114] <= wrong_col_114;
wrong_cnt[115] <= wrong_col_115;
wrong_cnt[116] <= wrong_col_116;
wrong_cnt[117] <= wrong_col_117;
wrong_cnt[118] <= wrong_col_118;
wrong_cnt[119] <= wrong_col_119;
wrong_cnt[120] <= wrong_col_120;
wrong_cnt[121] <= wrong_col_121;
wrong_cnt[122] <= wrong_col_122;
wrong_cnt[123] <= wrong_col_123;
wrong_cnt[124] <= wrong_col_124;
wrong_cnt[125] <= wrong_col_125;
wrong_cnt[126] <= wrong_col_126;
wrong_cnt[127] <= wrong_col_127;
wrong_cnt[128] <= wrong_col_128;
wrong_cnt[129] <= wrong_col_129;
wrong_cnt[130] <= wrong_col_130;
wrong_cnt[131] <= wrong_col_131;
wrong_cnt[132] <= wrong_col_132;
wrong_cnt[133] <= wrong_col_133;
wrong_cnt[134] <= wrong_col_134;
wrong_cnt[135] <= wrong_col_135;
wrong_cnt[136] <= wrong_col_136;
wrong_cnt[137] <= wrong_col_137;
wrong_cnt[138] <= wrong_col_138;
wrong_cnt[139] <= wrong_col_139;
wrong_cnt[140] <= wrong_col_140;
wrong_cnt[141] <= wrong_col_141;
wrong_cnt[142] <= wrong_col_142;
wrong_cnt[143] <= wrong_col_143;
wrong_cnt[144] <= wrong_col_144;
wrong_cnt[145] <= wrong_col_145;
wrong_cnt[146] <= wrong_col_146;
wrong_cnt[147] <= wrong_col_147;
wrong_cnt[148] <= wrong_col_148;
wrong_cnt[149] <= wrong_col_149;
wrong_cnt[150] <= wrong_col_150;
wrong_cnt[151] <= wrong_col_151;
wrong_cnt[152] <= wrong_col_152;
wrong_cnt[153] <= wrong_col_153;
wrong_cnt[154] <= wrong_col_154;
wrong_cnt[155] <= wrong_col_155;
wrong_cnt[156] <= wrong_col_156;
wrong_cnt[157] <= wrong_col_157;
wrong_cnt[158] <= wrong_col_158;
wrong_cnt[159] <= wrong_col_159;
wrong_cnt[160] <= wrong_col_160;
wrong_cnt[161] <= wrong_col_161;
wrong_cnt[162] <= wrong_col_162;
wrong_cnt[163] <= wrong_col_163;
wrong_cnt[164] <= wrong_col_164;
wrong_cnt[165] <= wrong_col_165;
wrong_cnt[166] <= wrong_col_166;
wrong_cnt[167] <= wrong_col_167;
wrong_cnt[168] <= wrong_col_168;
wrong_cnt[169] <= wrong_col_169;
wrong_cnt[170] <= wrong_col_170;
wrong_cnt[171] <= wrong_col_171;
wrong_cnt[172] <= wrong_col_172;
wrong_cnt[173] <= wrong_col_173;
wrong_cnt[174] <= wrong_col_174;
wrong_cnt[175] <= wrong_col_175;
wrong_cnt[176] <= wrong_col_176;
wrong_cnt[177] <= wrong_col_177;
wrong_cnt[178] <= wrong_col_178;
wrong_cnt[179] <= wrong_col_179;
wrong_cnt[180] <= wrong_col_180;
wrong_cnt[181] <= wrong_col_181;
wrong_cnt[182] <= wrong_col_182;
wrong_cnt[183] <= wrong_col_183;
wrong_cnt[184] <= wrong_col_184;
wrong_cnt[185] <= wrong_col_185;
wrong_cnt[186] <= wrong_col_186;
wrong_cnt[187] <= wrong_col_187;
wrong_cnt[188] <= wrong_col_188;
wrong_cnt[189] <= wrong_col_189;
wrong_cnt[190] <= wrong_col_190;
wrong_cnt[191] <= wrong_col_191;
wrong_cnt[192] <= wrong_col_192;
wrong_cnt[193] <= wrong_col_193;
wrong_cnt[194] <= wrong_col_194;
wrong_cnt[195] <= wrong_col_195;
wrong_cnt[196] <= wrong_col_196;
wrong_cnt[197] <= wrong_col_197;
wrong_cnt[198] <= wrong_col_198;
wrong_cnt[199] <= wrong_col_199;
wrong_cnt[200] <= wrong_col_200;
wrong_cnt[201] <= wrong_col_201;
wrong_cnt[202] <= wrong_col_202;
wrong_cnt[203] <= wrong_col_203;
wrong_cnt[204] <= wrong_col_204;
wrong_cnt[205] <= wrong_col_205;
wrong_cnt[206] <= wrong_col_206;
wrong_cnt[207] <= wrong_col_207;
wrong_cnt[208] <= wrong_col_208;
wrong_cnt[209] <= wrong_col_209;
wrong_cnt[210] <= wrong_col_210;
wrong_cnt[211] <= wrong_col_211;
wrong_cnt[212] <= wrong_col_212;
wrong_cnt[213] <= wrong_col_213;
wrong_cnt[214] <= wrong_col_214;
wrong_cnt[215] <= wrong_col_215;
wrong_cnt[216] <= wrong_col_216;
wrong_cnt[217] <= wrong_col_217;
wrong_cnt[218] <= wrong_col_218;
wrong_cnt[219] <= wrong_col_219;
wrong_cnt[220] <= wrong_col_220;
wrong_cnt[221] <= wrong_col_221;
wrong_cnt[222] <= wrong_col_222;
wrong_cnt[223] <= wrong_col_223;
wrong_cnt[224] <= wrong_col_224;
wrong_cnt[225] <= wrong_col_225;
wrong_cnt[226] <= wrong_col_226;
wrong_cnt[227] <= wrong_col_227;
wrong_cnt[228] <= wrong_col_228;
wrong_cnt[229] <= wrong_col_229;
wrong_cnt[230] <= wrong_col_230;
wrong_cnt[231] <= wrong_col_231;
wrong_cnt[232] <= wrong_col_232;
wrong_cnt[233] <= wrong_col_233;
wrong_cnt[234] <= wrong_col_234;
wrong_cnt[235] <= wrong_col_235;
wrong_cnt[236] <= wrong_col_236;
wrong_cnt[237] <= wrong_col_237;
wrong_cnt[238] <= wrong_col_238;
wrong_cnt[239] <= wrong_col_239;
wrong_cnt[240] <= wrong_col_240;
wrong_cnt[241] <= wrong_col_241;
wrong_cnt[242] <= wrong_col_242;
wrong_cnt[243] <= wrong_col_243;
wrong_cnt[244] <= wrong_col_244;
wrong_cnt[245] <= wrong_col_245;
wrong_cnt[246] <= wrong_col_246;
wrong_cnt[247] <= wrong_col_247;
wrong_cnt[248] <= wrong_col_248;
wrong_cnt[249] <= wrong_col_249;
wrong_cnt[250] <= wrong_col_250;
wrong_cnt[251] <= wrong_col_251;
wrong_cnt[252] <= wrong_col_252;
wrong_cnt[253] <= wrong_col_253;
wrong_cnt[254] <= wrong_col_254;
wrong_cnt[255] <= wrong_col_255;

state <= compare;

end


compare: begin
integer i;
for (i=0;i<256;i=i+1) begin
    if (wrong_cnt[i] >= check_cnt[i]) begin
        update_buffer[i] <= ~tx_buffer[i];
    end
    else begin
        update_buffer[i] <= tx_buffer[i];
    end
end
state <= update;

end


update: begin
integer i;
tx_buffer <= update_buffer;
iter_cnt <= iter_cnt + 1'b1;
if(iter_cnt >= iteration-2) begin
    valid_flag <= 1'b1;
    deout_reg <= tx_buffer;
    state <= decode;
end
else begin
    state <= getin;
end

end


decode: begin
valid_flag <= 1'b1;
deout_reg <= tx_buffer;
free_flag <= 1'b1;
iter_cnt <= 'd0;
iter_flag <= 1'b0;
state <= getin;

end

default: state <= init;

endcase


end //the end of biggest if
end //the end of always



endmodule

