module add_4(a1, a2, s);
input [2:0] a1, a2;
output wire [3:0] s;

assign s = a1 + a2;

endmodule
