module add_1.v(a1, a2, s);
input [0:0] a1, a2;
output wire [1:0] s;

assign s = a1 + a2;

endmodule
