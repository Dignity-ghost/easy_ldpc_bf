module add_16.v(a1, a2, s);
input [4:0] a1, a2;
output wire [5:0] s;

assign s = a1 + a2;

endmodule
